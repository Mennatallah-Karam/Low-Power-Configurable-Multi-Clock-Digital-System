module CLKBUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX20M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX14M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX16M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX1M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module DLY1X4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X1M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX12M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Thu Oct 24 02:39:05 2024
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN10_RST_N;
   wire FE_PHN9_RST_N;
   wire FE_PHN8_RST_N;
   wire FE_PHN4_scan_rst;
   wire FE_PHN3_scan_rst;
   wire FE_PHN0_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC10_RST_N (
	.Y(FE_PHN10_RST_N),
	.A(FE_PHN9_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC9_RST_N (
	.Y(FE_PHN9_RST_N),
	.A(FE_PHN8_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC8_RST_N (
	.Y(FE_PHN8_RST_N),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC4_scan_rst (
	.Y(FE_PHN4_scan_rst),
	.A(FE_PHN3_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC3_scan_rst (
	.Y(FE_PHN3_scan_rst),
	.A(FE_PHN0_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_scan_rst (
	.Y(FE_PHN0_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN4_scan_rst),
	.A(FE_PHN10_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_scan_rst;
   wire FE_PHN6_scan_rst;
   wire FE_PHN2_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC7_scan_rst (
	.Y(FE_PHN7_scan_rst),
	.A(FE_PHN6_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC6_scan_rst (
	.Y(FE_PHN6_scan_rst),
	.A(FE_PHN2_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_scan_rst (
	.Y(FE_PHN2_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X6M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN7_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN5_scan_rst;
   wire FE_PHN1_scan_rst;
   wire N0;

   assign N0 = SEL ;

   // Module instantiations
   DLY4X1M FE_PHC5_scan_rst (
	.Y(FE_PHN5_scan_rst),
	.A(FE_PHN1_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC1_scan_rst (
	.Y(FE_PHN1_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(N0),
	.B(FE_PHN5_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_0 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \FFs[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FFs_reg[1]  (
	.SI(\FFs[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\FFs[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FFs_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\FFs[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYNC_test_1 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_se, 
	UART_SCAN_CLK__L3_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   input test_se;
   input UART_SCAN_CLK__L3_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \FFs[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FFs_reg[1]  (
	.SI(\FFs[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\FFs[0] ),
	.CK(UART_SCAN_CLK__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \FFs_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\FFs[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DataSynchronizer_BUS_WIDTH8_test_1 (
	Unsync_bus, 
	bus_enable, 
	CLK, 
	RST, 
	sync_bus, 
	enable_pulse, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN2_SYNC_SCAN_RST1, 
	VDD, 
	VSS);
   input [7:0] Unsync_bus;
   input bus_enable;
   input CLK;
   input RST;
   output [7:0] sync_bus;
   output enable_pulse;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN2_SYNC_SCAN_RST1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN12_n20__Exclude_0_NET;
   wire sync_enable_F3;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire [1:0] sync_enable_FF;

   assign test_so = sync_enable_FF[1] ;

   // Module instantiations
   DLY4X1M FE_PHC12_n20__Exclude_0_NET (
	.Y(FE_PHN12_n20__Exclude_0_NET),
	.A(test_si), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n10),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U4 (
	.Y(n1),
	.B(sync_enable_FF[1]),
	.AN(sync_enable_F3), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U5 (
	.Y(n2),
	.B1(n1),
	.B0(sync_bus[0]),
	.A1(n10),
	.A0(Unsync_bus[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n3),
	.B1(n1),
	.B0(sync_bus[1]),
	.A1(n10),
	.A0(Unsync_bus[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n4),
	.B1(n1),
	.B0(sync_bus[2]),
	.A1(n10),
	.A0(Unsync_bus[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n5),
	.B1(n1),
	.B0(sync_bus[3]),
	.A1(n10),
	.A0(Unsync_bus[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n6),
	.B1(n1),
	.B0(sync_bus[4]),
	.A1(n10),
	.A0(Unsync_bus[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n7),
	.B1(n1),
	.B0(sync_bus[5]),
	.A1(n10),
	.A0(Unsync_bus[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n8),
	.B1(n1),
	.B0(sync_bus[6]),
	.A1(n10),
	.A0(Unsync_bus[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n9),
	.B1(n1),
	.B0(sync_bus[7]),
	.A1(n10),
	.A0(Unsync_bus[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sync_enable_F3_reg (
	.SI(sync_bus[7]),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(sync_enable_F3),
	.D(sync_enable_FF[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_enable_FF_reg[1]  (
	.SI(sync_enable_FF[0]),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(sync_enable_FF[1]),
	.D(sync_enable_FF[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[7]  (
	.SI(sync_bus[6]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[7]),
	.D(n9),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[4]  (
	.SI(sync_bus[3]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[4]),
	.D(n6),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[6]  (
	.SI(sync_bus[5]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[6]),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[5]  (
	.SI(sync_bus[4]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[5]),
	.D(n7),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[3]  (
	.SI(sync_bus[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[3]),
	.D(n5),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[2]  (
	.SI(sync_bus[1]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_bus[2]),
	.D(n4),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[0]  (
	.SI(enable_pulse),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(sync_bus[0]),
	.D(n2),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[1]  (
	.SI(sync_bus[0]),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(sync_bus[1]),
	.D(n3),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_pulse_reg (
	.SI(FE_PHN12_n20__Exclude_0_NET),
	.SE(test_se),
	.RN(RST),
	.Q(enable_pulse),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_enable_FF_reg[0]  (
	.SI(sync_enable_F3),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(sync_enable_FF[0]),
	.D(bus_enable),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_TOP_DATA_WIDTH8_test_1 (
	wclk, 
	rclk, 
	wrst_n, 
	rrst_n, 
	winc, 
	rinc, 
	wdata, 
	rdata, 
	wfull, 
	empty, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN2_SYNC_SCAN_RST1, 
	REF_SCAN_CLK__L6_N11, 
	REF_SCAN_CLK__L6_N12, 
	REF_SCAN_CLK__L6_N13, 
	REF_SCAN_CLK__L6_N4, 
	REF_SCAN_CLK__L6_N5, 
	REF_SCAN_CLK__L6_N6, 
	VDD, 
	VSS);
   input wclk;
   input rclk;
   input wrst_n;
   input rrst_n;
   input winc;
   input rinc;
   input [7:0] wdata;
   output [7:0] rdata;
   output wfull;
   output empty;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN2_SYNC_SCAN_RST1;
   input REF_SCAN_CLK__L6_N11;
   input REF_SCAN_CLK__L6_N12;
   input REF_SCAN_CLK__L6_N13;
   input REF_SCAN_CLK__L6_N4;
   input REF_SCAN_CLK__L6_N5;
   input REF_SCAN_CLK__L6_N6;
   inout VDD;
   inout VSS;

   // Internal wires
   wire wclken;
   wire n3;
   wire [3:0] sync_r2w;
   wire [3:0] wptr_gray;
   wire [2:0] waddr;
   wire [3:0] sync_w2r;
   wire [2:0] raddr;
   wire [3:0] rptr_gray;

   assign test_so2 = sync_w2r[3] ;

   // Module instantiations
   FIFO_WR_FIFO_DEPTH8_ADDR_WIDTH4_test_1 fifo_wr (
	.wdata({ wdata[7],
		wdata[6],
		wdata[5],
		wdata[4],
		wdata[3],
		wdata[2],
		wdata[1],
		wdata[0] }),
	.wclk(REF_SCAN_CLK__L6_N12),
	.wrst_n(FE_OFN2_SYNC_SCAN_RST1),
	.winc(winc),
	.rptr_gray({ sync_r2w[3],
		sync_r2w[2],
		sync_r2w[1],
		sync_r2w[0] }),
	.wptr_gray({ wptr_gray[3],
		wptr_gray[2],
		wptr_gray[1],
		wptr_gray[0] }),
	.waddr({ waddr[2],
		waddr[1],
		waddr[0] }),
	.wclken(wclken),
	.wfull(wfull),
	.test_si(rptr_gray[3]),
	.test_se(test_se),
	.REF_SCAN_CLK__L6_N13(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_RD_FIFO_DEPTH8_ADDR_WIDTH4_test_1 fifo_rd (
	.wptr_gray({ sync_w2r[3],
		sync_w2r[2],
		sync_w2r[1],
		sync_w2r[0] }),
	.rclk(rclk),
	.rrst_n(rrst_n),
	.rinc(rinc),
	.raddr({ raddr[2],
		raddr[1],
		raddr[0] }),
	.rptr_gray({ rptr_gray[3],
		rptr_gray[2],
		rptr_gray[1],
		rptr_gray[0] }),
	.empty(empty),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_SYNC_WIDTH4_test_0 sync_rptr_gray_to_wptr_gray (
	.RST(FE_OFN2_SYNC_SCAN_RST1),
	.CLK(REF_SCAN_CLK__L6_N13),
	.async_signal({ rptr_gray[3],
		rptr_gray[2],
		rptr_gray[1],
		rptr_gray[0] }),
	.sync_signal({ sync_r2w[3],
		sync_r2w[2],
		sync_r2w[1],
		sync_r2w[0] }),
	.test_si(wptr_gray[3]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_SYNC_WIDTH4_test_1 sync_wptr_gray_to_rptr_gray (
	.RST(rrst_n),
	.CLK(rclk),
	.async_signal({ wptr_gray[3],
		wptr_gray[2],
		wptr_gray[1],
		wptr_gray[0] }),
	.sync_signal({ sync_w2r[3],
		sync_w2r[2],
		sync_w2r[1],
		sync_w2r[0] }),
	.test_si(sync_r2w[3]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_MEM_CNTRL_DATA_WIDTH8_FIFO_DEPTH8_ADDR_WIDTH4_test_1 fifo_mem (
	.wdata({ wdata[7],
		wdata[6],
		wdata[5],
		wdata[4],
		wdata[3],
		wdata[2],
		wdata[1],
		wdata[0] }),
	.waddr({ waddr[2],
		waddr[1],
		waddr[0] }),
	.raddr({ raddr[2],
		raddr[1],
		raddr[0] }),
	.wclk(wclk),
	.rclk(rclk),
	.wrst_n(wrst_n),
	.wclken(wclken),
	.rdata({ rdata[7],
		rdata[6],
		rdata[5],
		rdata[4],
		rdata[3],
		rdata[2],
		rdata[1],
		rdata[0] }),
	.test_si2(test_si2),
	.test_si1(test_si1),
	.test_so2(n3),
	.test_so1(test_so1),
	.test_se(test_se),
	.FE_OFN2_SYNC_SCAN_RST1(FE_OFN2_SYNC_SCAN_RST1),
	.REF_SCAN_CLK__L6_N11(REF_SCAN_CLK__L6_N11),
	.REF_SCAN_CLK__L6_N12(REF_SCAN_CLK__L6_N12),
	.REF_SCAN_CLK__L6_N13(REF_SCAN_CLK__L6_N13),
	.REF_SCAN_CLK__L6_N4(REF_SCAN_CLK__L6_N4),
	.REF_SCAN_CLK__L6_N5(REF_SCAN_CLK__L6_N5),
	.REF_SCAN_CLK__L6_N6(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_WR_FIFO_DEPTH8_ADDR_WIDTH4_test_1 (
	wdata, 
	wclk, 
	wrst_n, 
	winc, 
	rptr_gray, 
	wptr_gray, 
	waddr, 
	wclken, 
	wfull, 
	test_si, 
	test_se, 
	REF_SCAN_CLK__L6_N13, 
	VDD, 
	VSS);
   input [7:0] wdata;
   input wclk;
   input wrst_n;
   input winc;
   input [3:0] rptr_gray;
   output [3:0] wptr_gray;
   output [2:0] waddr;
   output wclken;
   output wfull;
   input test_si;
   input test_se;
   input REF_SCAN_CLK__L6_N13;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;

   // Module instantiations
   INVX2M U3 (
	.Y(wclken),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U4 (
	.Y(n3),
	.B(n2),
	.A(winc), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(wfull),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(n7),
	.B(rptr_gray[1]),
	.A(wptr_gray[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(wptr_gray[0]),
	.B(waddr[1]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U8 (
	.Y(n6),
	.B(n1),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n12),
	.B(n5),
	.A(waddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n11),
	.B(n4),
	.A(wptr_gray[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U11 (
	.Y(n4),
	.B(waddr[2]),
	.AN(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U12 (
	.Y(n2),
	.D(n10),
	.C(n9),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(n10),
	.B(rptr_gray[3]),
	.A(wptr_gray[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U14 (
	.Y(n8),
	.B(rptr_gray[0]),
	.A(wptr_gray[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(n9),
	.B(wptr_gray[2]),
	.A(rptr_gray[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(n5),
	.B(waddr[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(wptr_gray[2]),
	.B(waddr[2]),
	.A(wptr_gray[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(wptr_gray[1]),
	.B(waddr[2]),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(n13),
	.B(n6),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U20 (
	.Y(n14),
	.B(n3),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg[3]  (
	.SI(waddr[2]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(wptr_gray[3]),
	.D(n11),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg[2]  (
	.SI(waddr[1]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(waddr[2]),
	.D(n12),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \wptr_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(wrst_n),
	.QN(n1),
	.Q(waddr[0]),
	.D(n14),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wptr_reg[1]  (
	.SI(waddr[0]),
	.SE(test_se),
	.RN(wrst_n),
	.Q(waddr[1]),
	.D(n13),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_RD_FIFO_DEPTH8_ADDR_WIDTH4_test_1 (
	wptr_gray, 
	rclk, 
	rrst_n, 
	rinc, 
	raddr, 
	rptr_gray, 
	empty, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [3:0] wptr_gray;
   input rclk;
   input rrst_n;
   input rinc;
   output [2:0] raddr;
   output [3:0] rptr_gray;
   output empty;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;

   // Module instantiations
   XNOR2X2M U4 (
	.Y(n7),
	.B(wptr_gray[1]),
	.A(rptr_gray[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(rptr_gray[0]),
	.B(raddr[1]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n4),
	.B(n1),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n11),
	.B(n2),
	.A(rptr_gray[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U8 (
	.Y(n2),
	.B(raddr[2]),
	.AN(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U9 (
	.Y(empty),
	.D(n10),
	.C(n9),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n9),
	.B(wptr_gray[3]),
	.A(rptr_gray[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U11 (
	.Y(n10),
	.B(wptr_gray[2]),
	.A(rptr_gray[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U12 (
	.Y(n8),
	.B(wptr_gray[0]),
	.A(rptr_gray[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U13 (
	.Y(n3),
	.B(raddr[1]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(n5),
	.B(empty),
	.A(rinc), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(rptr_gray[1]),
	.B(raddr[2]),
	.A(raddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(rptr_gray[2]),
	.B(raddr[2]),
	.A(rptr_gray[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U17 (
	.Y(n12),
	.B(n3),
	.A(raddr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(n13),
	.B(n4),
	.A(raddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(n14),
	.B(n5),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rptr_reg[3]  (
	.SI(raddr[2]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(rptr_gray[3]),
	.D(n11),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \rptr_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rrst_n),
	.QN(n1),
	.Q(raddr[0]),
	.D(n14),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rptr_reg[2]  (
	.SI(raddr[1]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddr[2]),
	.D(n12),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \rptr_reg[1]  (
	.SI(raddr[0]),
	.SE(test_se),
	.RN(rrst_n),
	.Q(raddr[1]),
	.D(n13),
	.CK(rclk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_SYNC_WIDTH4_test_0 (
	RST, 
	CLK, 
	async_signal, 
	sync_signal, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   input [3:0] async_signal;
   output [3:0] sync_signal;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [3:0] sync_ff1;

   // Module instantiations
   SDFFRQX2M \sync_ff2_reg[1]  (
	.SI(sync_signal[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[1]),
	.D(sync_ff1[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff2_reg[0]  (
	.SI(sync_ff1[3]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[0]),
	.D(sync_ff1[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff2_reg[2]  (
	.SI(sync_signal[1]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[2]),
	.D(sync_ff1[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff2_reg[3]  (
	.SI(sync_signal[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[3]),
	.D(sync_ff1[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[3]  (
	.SI(sync_ff1[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[3]),
	.D(async_signal[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[2]  (
	.SI(sync_ff1[1]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[2]),
	.D(async_signal[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[1]  (
	.SI(sync_ff1[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[1]),
	.D(async_signal[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[0]),
	.D(async_signal[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_SYNC_WIDTH4_test_1 (
	RST, 
	CLK, 
	async_signal, 
	sync_signal, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   input [3:0] async_signal;
   output [3:0] sync_signal;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [3:0] sync_ff1;

   // Module instantiations
   SDFFRQX2M \sync_ff2_reg[3]  (
	.SI(sync_signal[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[3]),
	.D(sync_ff1[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff2_reg[2]  (
	.SI(sync_signal[1]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[2]),
	.D(sync_ff1[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff2_reg[1]  (
	.SI(sync_signal[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[1]),
	.D(sync_ff1[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff2_reg[0]  (
	.SI(sync_ff1[3]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_signal[0]),
	.D(sync_ff1[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[3]  (
	.SI(sync_ff1[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[3]),
	.D(async_signal[3]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[2]  (
	.SI(sync_ff1[1]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[2]),
	.D(async_signal[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[1]  (
	.SI(sync_ff1[0]),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[1]),
	.D(async_signal[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_ff1_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(sync_ff1[0]),
	.D(async_signal[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_MEM_CNTRL_DATA_WIDTH8_FIFO_DEPTH8_ADDR_WIDTH4_test_1 (
	wdata, 
	waddr, 
	raddr, 
	wclk, 
	rclk, 
	wrst_n, 
	wclken, 
	rdata, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN2_SYNC_SCAN_RST1, 
	REF_SCAN_CLK__L6_N11, 
	REF_SCAN_CLK__L6_N12, 
	REF_SCAN_CLK__L6_N13, 
	REF_SCAN_CLK__L6_N4, 
	REF_SCAN_CLK__L6_N5, 
	REF_SCAN_CLK__L6_N6, 
	VDD, 
	VSS);
   input [7:0] wdata;
   input [2:0] waddr;
   input [2:0] raddr;
   input wclk;
   input rclk;
   input wrst_n;
   input wclken;
   output [7:0] rdata;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN2_SYNC_SCAN_RST1;
   input REF_SCAN_CLK__L6_N11;
   input REF_SCAN_CLK__L6_N12;
   input REF_SCAN_CLK__L6_N13;
   input REF_SCAN_CLK__L6_N4;
   input REF_SCAN_CLK__L6_N5;
   input REF_SCAN_CLK__L6_N6;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN7_SO_3_;
   wire N10;
   wire N11;
   wire N12;
   wire \fifo_mem[0][7] ;
   wire \fifo_mem[0][6] ;
   wire \fifo_mem[0][5] ;
   wire \fifo_mem[0][4] ;
   wire \fifo_mem[0][3] ;
   wire \fifo_mem[0][2] ;
   wire \fifo_mem[0][1] ;
   wire \fifo_mem[0][0] ;
   wire \fifo_mem[1][7] ;
   wire \fifo_mem[1][6] ;
   wire \fifo_mem[1][5] ;
   wire \fifo_mem[1][4] ;
   wire \fifo_mem[1][3] ;
   wire \fifo_mem[1][2] ;
   wire \fifo_mem[1][1] ;
   wire \fifo_mem[1][0] ;
   wire \fifo_mem[2][7] ;
   wire \fifo_mem[2][6] ;
   wire \fifo_mem[2][5] ;
   wire \fifo_mem[2][4] ;
   wire \fifo_mem[2][3] ;
   wire \fifo_mem[2][2] ;
   wire \fifo_mem[2][1] ;
   wire \fifo_mem[2][0] ;
   wire \fifo_mem[3][7] ;
   wire \fifo_mem[3][6] ;
   wire \fifo_mem[3][5] ;
   wire \fifo_mem[3][4] ;
   wire \fifo_mem[3][3] ;
   wire \fifo_mem[3][2] ;
   wire \fifo_mem[3][1] ;
   wire \fifo_mem[3][0] ;
   wire \fifo_mem[4][7] ;
   wire \fifo_mem[4][6] ;
   wire \fifo_mem[4][5] ;
   wire \fifo_mem[4][4] ;
   wire \fifo_mem[4][3] ;
   wire \fifo_mem[4][2] ;
   wire \fifo_mem[4][1] ;
   wire \fifo_mem[4][0] ;
   wire \fifo_mem[5][7] ;
   wire \fifo_mem[5][6] ;
   wire \fifo_mem[5][5] ;
   wire \fifo_mem[5][4] ;
   wire \fifo_mem[5][3] ;
   wire \fifo_mem[5][2] ;
   wire \fifo_mem[5][1] ;
   wire \fifo_mem[5][0] ;
   wire \fifo_mem[6][7] ;
   wire \fifo_mem[6][6] ;
   wire \fifo_mem[6][5] ;
   wire \fifo_mem[6][4] ;
   wire \fifo_mem[6][3] ;
   wire \fifo_mem[6][2] ;
   wire \fifo_mem[6][1] ;
   wire \fifo_mem[6][0] ;
   wire \fifo_mem[7][7] ;
   wire \fifo_mem[7][6] ;
   wire \fifo_mem[7][5] ;
   wire \fifo_mem[7][4] ;
   wire \fifo_mem[7][3] ;
   wire \fifo_mem[7][2] ;
   wire \fifo_mem[7][1] ;
   wire \fifo_mem[7][0] ;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;

   assign N10 = raddr[0] ;
   assign N11 = raddr[1] ;
   assign N12 = raddr[2] ;
   assign test_so1 = \fifo_mem[4][4]  ;
   assign test_so2 = \fifo_mem[7][7]  ;

   // Module instantiations
   BUFX10M FE_OFC7_SO_3_ (
	.Y(\fifo_mem[4][4] ),
	.A(FE_OFN7_SO_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U14 (
	.Y(n15),
	.C(n12),
	.B(n106),
	.A(n105), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U15 (
	.Y(n20),
	.C(n17),
	.B(n106),
	.A(n105), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U16 (
	.Y(n17),
	.B(waddr[2]),
	.AN(wclken), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U17 (
	.Y(n77),
	.B1(n20),
	.B0(n114),
	.A1N(n20),
	.A0N(\fifo_mem[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U18 (
	.Y(n78),
	.B1(n20),
	.B0(n113),
	.A1N(n20),
	.A0N(\fifo_mem[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U19 (
	.Y(n79),
	.B1(n20),
	.B0(n112),
	.A1N(n20),
	.A0N(\fifo_mem[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U20 (
	.Y(n80),
	.B1(n20),
	.B0(n111),
	.A1N(n20),
	.A0N(\fifo_mem[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U21 (
	.Y(n81),
	.B1(n20),
	.B0(n110),
	.A1N(n20),
	.A0N(\fifo_mem[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U22 (
	.Y(n82),
	.B1(n20),
	.B0(n109),
	.A1N(n20),
	.A0N(\fifo_mem[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U23 (
	.Y(n83),
	.B1(n20),
	.B0(n108),
	.A1N(n20),
	.A0N(\fifo_mem[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U24 (
	.Y(n84),
	.B1(n20),
	.B0(n107),
	.A1N(n20),
	.A0N(\fifo_mem[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U25 (
	.Y(n45),
	.B1(n15),
	.B0(n114),
	.A1N(n15),
	.A0N(\fifo_mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U26 (
	.Y(n46),
	.B1(n15),
	.B0(n113),
	.A1N(n15),
	.A0N(\fifo_mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U27 (
	.Y(n47),
	.B1(n15),
	.B0(n112),
	.A1N(n15),
	.A0N(\fifo_mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U28 (
	.Y(n48),
	.B1(n15),
	.B0(n111),
	.A1N(n15),
	.A0N(\fifo_mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U29 (
	.Y(n49),
	.B1(n15),
	.B0(n110),
	.A1N(n15),
	.A0N(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U30 (
	.Y(n50),
	.B1(n15),
	.B0(n109),
	.A1N(n15),
	.A0N(\fifo_mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U31 (
	.Y(n51),
	.B1(n15),
	.B0(n108),
	.A1N(n15),
	.A0N(\fifo_mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U32 (
	.Y(n52),
	.B1(n15),
	.B0(n107),
	.A1N(n15),
	.A0N(\fifo_mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U33 (
	.Y(n91),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n114),
	.A(wdata[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U35 (
	.Y(n113),
	.A(wdata[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n112),
	.A(wdata[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n111),
	.A(wdata[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n110),
	.A(wdata[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n109),
	.A(wdata[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n108),
	.A(wdata[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n107),
	.A(wdata[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U43 (
	.Y(n19),
	.C(n17),
	.B(n106),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U44 (
	.Y(n29),
	.B1(n13),
	.B0(n114),
	.A1N(n13),
	.A0N(\fifo_mem[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U45 (
	.Y(n30),
	.B1(n13),
	.B0(n113),
	.A1N(n13),
	.A0N(\fifo_mem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U46 (
	.Y(n31),
	.B1(n13),
	.B0(n112),
	.A1N(n13),
	.A0N(\fifo_mem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U47 (
	.Y(n32),
	.B1(n13),
	.B0(n111),
	.A1N(n13),
	.A0N(\fifo_mem[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U48 (
	.Y(n33),
	.B1(n13),
	.B0(n110),
	.A1N(n13),
	.A0N(\fifo_mem[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U49 (
	.Y(n34),
	.B1(n13),
	.B0(n109),
	.A1N(n13),
	.A0N(\fifo_mem[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U50 (
	.Y(n35),
	.B1(n13),
	.B0(n108),
	.A1N(n13),
	.A0N(\fifo_mem[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U51 (
	.Y(n36),
	.B1(n13),
	.B0(n107),
	.A1N(n13),
	.A0N(\fifo_mem[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U52 (
	.Y(n37),
	.B1(n14),
	.B0(n114),
	.A1N(n14),
	.A0N(\fifo_mem[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U53 (
	.Y(n38),
	.B1(n14),
	.B0(n113),
	.A1N(n14),
	.A0N(\fifo_mem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U54 (
	.Y(n39),
	.B1(n14),
	.B0(n112),
	.A1N(n14),
	.A0N(\fifo_mem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U55 (
	.Y(n40),
	.B1(n14),
	.B0(n111),
	.A1N(n14),
	.A0N(\fifo_mem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U56 (
	.Y(n41),
	.B1(n14),
	.B0(n110),
	.A1N(n14),
	.A0N(\fifo_mem[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U57 (
	.Y(n42),
	.B1(n14),
	.B0(n109),
	.A1N(n14),
	.A0N(\fifo_mem[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U58 (
	.Y(n43),
	.B1(n14),
	.B0(n108),
	.A1N(n14),
	.A0N(\fifo_mem[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U59 (
	.Y(n44),
	.B1(n14),
	.B0(n107),
	.A1N(n14),
	.A0N(\fifo_mem[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U60 (
	.Y(n53),
	.B1(n16),
	.B0(n114),
	.A1N(n16),
	.A0N(\fifo_mem[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U61 (
	.Y(n54),
	.B1(n16),
	.B0(n113),
	.A1N(n16),
	.A0N(\fifo_mem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U62 (
	.Y(n55),
	.B1(n16),
	.B0(n112),
	.A1N(n16),
	.A0N(\fifo_mem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U63 (
	.Y(n56),
	.B1(n16),
	.B0(n111),
	.A1N(n16),
	.A0N(\fifo_mem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U64 (
	.Y(n57),
	.B1(n16),
	.B0(n110),
	.A1N(n16),
	.A0N(\fifo_mem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U65 (
	.Y(n58),
	.B1(n16),
	.B0(n109),
	.A1N(n16),
	.A0N(\fifo_mem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U66 (
	.Y(n59),
	.B1(n16),
	.B0(n108),
	.A1N(n16),
	.A0N(\fifo_mem[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U67 (
	.Y(n60),
	.B1(n16),
	.B0(n107),
	.A1N(n16),
	.A0N(\fifo_mem[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U68 (
	.Y(n61),
	.B1(n18),
	.B0(n114),
	.A1N(n18),
	.A0N(\fifo_mem[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U69 (
	.Y(n62),
	.B1(n18),
	.B0(n113),
	.A1N(n18),
	.A0N(\fifo_mem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U70 (
	.Y(n63),
	.B1(n18),
	.B0(n112),
	.A1N(n18),
	.A0N(\fifo_mem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U71 (
	.Y(n64),
	.B1(n18),
	.B0(n111),
	.A1N(n18),
	.A0N(\fifo_mem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U72 (
	.Y(n65),
	.B1(n18),
	.B0(n110),
	.A1N(n18),
	.A0N(\fifo_mem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U73 (
	.Y(n66),
	.B1(n18),
	.B0(n109),
	.A1N(n18),
	.A0N(\fifo_mem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U74 (
	.Y(n67),
	.B1(n18),
	.B0(n108),
	.A1N(n18),
	.A0N(\fifo_mem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U75 (
	.Y(n68),
	.B1(n18),
	.B0(n107),
	.A1N(n18),
	.A0N(\fifo_mem[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U76 (
	.Y(n69),
	.B1(n19),
	.B0(n114),
	.A1N(n19),
	.A0N(\fifo_mem[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U77 (
	.Y(n70),
	.B1(n19),
	.B0(n113),
	.A1N(n19),
	.A0N(\fifo_mem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U78 (
	.Y(n71),
	.B1(n19),
	.B0(n112),
	.A1N(n19),
	.A0N(\fifo_mem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U79 (
	.Y(n72),
	.B1(n19),
	.B0(n111),
	.A1N(n19),
	.A0N(\fifo_mem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U80 (
	.Y(n73),
	.B1(n19),
	.B0(n110),
	.A1N(n19),
	.A0N(\fifo_mem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U81 (
	.Y(n74),
	.B1(n19),
	.B0(n109),
	.A1N(n19),
	.A0N(\fifo_mem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U82 (
	.Y(n75),
	.B1(n19),
	.B0(n108),
	.A1N(n19),
	.A0N(\fifo_mem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U83 (
	.Y(n76),
	.B1(n19),
	.B0(n107),
	.A1N(n19),
	.A0N(\fifo_mem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n21),
	.B1(n114),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n22),
	.B1(n113),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n23),
	.B1(n112),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n24),
	.B1(n111),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n25),
	.B1(n110),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n26),
	.B1(n109),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n27),
	.B1(n108),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n28),
	.B1(n107),
	.B0(n11),
	.A1N(n11),
	.A0N(\fifo_mem[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U92 (
	.Y(n12),
	.B(waddr[2]),
	.A(wclken), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U93 (
	.Y(n14),
	.C(waddr[0]),
	.B(n106),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U94 (
	.Y(n13),
	.C(waddr[1]),
	.B(n105),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U95 (
	.Y(n16),
	.C(n17),
	.B(waddr[0]),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U96 (
	.Y(n18),
	.C(n17),
	.B(n105),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U97 (
	.Y(n11),
	.C(waddr[1]),
	.B(n12),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U98 (
	.Y(rdata[0]),
	.S0(N12),
	.B(n1),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U99 (
	.Y(n2),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][0] ),
	.C(\fifo_mem[2][0] ),
	.B(\fifo_mem[1][0] ),
	.A(\fifo_mem[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U100 (
	.Y(n1),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][0] ),
	.C(\fifo_mem[6][0] ),
	.B(\fifo_mem[5][0] ),
	.A(\fifo_mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U101 (
	.Y(rdata[1]),
	.S0(N12),
	.B(n3),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U102 (
	.Y(n4),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][1] ),
	.C(\fifo_mem[2][1] ),
	.B(\fifo_mem[1][1] ),
	.A(\fifo_mem[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U103 (
	.Y(n3),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][1] ),
	.C(\fifo_mem[6][1] ),
	.B(\fifo_mem[5][1] ),
	.A(\fifo_mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U104 (
	.Y(rdata[2]),
	.S0(N12),
	.B(n5),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U105 (
	.Y(n6),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][2] ),
	.C(\fifo_mem[2][2] ),
	.B(\fifo_mem[1][2] ),
	.A(\fifo_mem[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U106 (
	.Y(n5),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][2] ),
	.C(\fifo_mem[6][2] ),
	.B(\fifo_mem[5][2] ),
	.A(\fifo_mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U107 (
	.Y(rdata[3]),
	.S0(N12),
	.B(n7),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U108 (
	.Y(n8),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][3] ),
	.C(\fifo_mem[2][3] ),
	.B(\fifo_mem[1][3] ),
	.A(\fifo_mem[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U109 (
	.Y(n7),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][3] ),
	.C(\fifo_mem[6][3] ),
	.B(\fifo_mem[5][3] ),
	.A(\fifo_mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U110 (
	.Y(rdata[4]),
	.S0(N12),
	.B(n9),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U111 (
	.Y(n10),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][4] ),
	.C(\fifo_mem[2][4] ),
	.B(\fifo_mem[1][4] ),
	.A(\fifo_mem[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U112 (
	.Y(n9),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][4] ),
	.C(\fifo_mem[6][4] ),
	.B(\fifo_mem[5][4] ),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U113 (
	.Y(rdata[5]),
	.S0(N12),
	.B(n85),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U114 (
	.Y(n86),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][5] ),
	.C(\fifo_mem[2][5] ),
	.B(\fifo_mem[1][5] ),
	.A(\fifo_mem[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U115 (
	.Y(n85),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][5] ),
	.C(\fifo_mem[6][5] ),
	.B(\fifo_mem[5][5] ),
	.A(\fifo_mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U116 (
	.Y(rdata[6]),
	.S0(N12),
	.B(n87),
	.A(n88), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U117 (
	.Y(n88),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][6] ),
	.C(\fifo_mem[2][6] ),
	.B(\fifo_mem[1][6] ),
	.A(\fifo_mem[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U118 (
	.Y(n87),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][6] ),
	.C(\fifo_mem[6][6] ),
	.B(\fifo_mem[5][6] ),
	.A(\fifo_mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U119 (
	.Y(rdata[7]),
	.S0(N12),
	.B(n89),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U120 (
	.Y(n90),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[3][7] ),
	.C(\fifo_mem[2][7] ),
	.B(\fifo_mem[1][7] ),
	.A(\fifo_mem[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U121 (
	.Y(n89),
	.S1(N11),
	.S0(n91),
	.D(\fifo_mem[7][7] ),
	.C(\fifo_mem[6][7] ),
	.B(\fifo_mem[5][7] ),
	.A(\fifo_mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U122 (
	.Y(n105),
	.A(waddr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U123 (
	.Y(n106),
	.A(waddr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][7]  (
	.SI(\fifo_mem[1][6] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][7] ),
	.D(n76),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][6]  (
	.SI(\fifo_mem[1][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][6] ),
	.D(n75),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][5]  (
	.SI(\fifo_mem[1][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][5] ),
	.D(n74),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][4]  (
	.SI(\fifo_mem[1][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][4] ),
	.D(n73),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][3]  (
	.SI(\fifo_mem[1][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][3] ),
	.D(n72),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][2]  (
	.SI(\fifo_mem[1][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][2] ),
	.D(n71),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][1]  (
	.SI(\fifo_mem[1][0] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[1][1] ),
	.D(n70),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[1][0]  (
	.SI(\fifo_mem[0][7] ),
	.SE(n122),
	.RN(wrst_n),
	.Q(\fifo_mem[1][0] ),
	.D(n69),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][7]  (
	.SI(\fifo_mem[5][6] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[5][7] ),
	.D(n44),
	.CK(REF_SCAN_CLK__L6_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][6]  (
	.SI(\fifo_mem[5][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[5][6] ),
	.D(n43),
	.CK(REF_SCAN_CLK__L6_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][5]  (
	.SI(\fifo_mem[5][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[5][5] ),
	.D(n42),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][4]  (
	.SI(\fifo_mem[5][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[5][4] ),
	.D(n41),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][3]  (
	.SI(\fifo_mem[5][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[5][3] ),
	.D(n40),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][2]  (
	.SI(\fifo_mem[5][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[5][2] ),
	.D(n39),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][1]  (
	.SI(\fifo_mem[5][0] ),
	.SE(n119),
	.RN(wrst_n),
	.Q(\fifo_mem[5][1] ),
	.D(n38),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[5][0]  (
	.SI(\fifo_mem[4][7] ),
	.SE(n122),
	.RN(wrst_n),
	.Q(\fifo_mem[5][0] ),
	.D(n37),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][7]  (
	.SI(\fifo_mem[3][6] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][7] ),
	.D(n60),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][6]  (
	.SI(\fifo_mem[3][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][6] ),
	.D(n59),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][5]  (
	.SI(\fifo_mem[3][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][5] ),
	.D(n58),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][4]  (
	.SI(\fifo_mem[3][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][4] ),
	.D(n57),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][3]  (
	.SI(\fifo_mem[3][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][3] ),
	.D(n56),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][2]  (
	.SI(\fifo_mem[3][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][2] ),
	.D(n55),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][1]  (
	.SI(\fifo_mem[3][0] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][1] ),
	.D(n54),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[3][0]  (
	.SI(\fifo_mem[2][7] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[3][0] ),
	.D(n53),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][7]  (
	.SI(\fifo_mem[7][6] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[7][7] ),
	.D(n28),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][6]  (
	.SI(\fifo_mem[7][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[7][6] ),
	.D(n27),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][5]  (
	.SI(\fifo_mem[7][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[7][5] ),
	.D(n26),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][4]  (
	.SI(\fifo_mem[7][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[7][4] ),
	.D(n25),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][3]  (
	.SI(\fifo_mem[7][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[7][3] ),
	.D(n24),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][2]  (
	.SI(\fifo_mem[7][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[7][2] ),
	.D(n23),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][1]  (
	.SI(\fifo_mem[7][0] ),
	.SE(n119),
	.RN(wrst_n),
	.Q(\fifo_mem[7][1] ),
	.D(n22),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[7][0]  (
	.SI(\fifo_mem[6][7] ),
	.SE(n122),
	.RN(wrst_n),
	.Q(\fifo_mem[7][0] ),
	.D(n21),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][7]  (
	.SI(\fifo_mem[2][6] ),
	.SE(n121),
	.RN(wrst_n),
	.Q(\fifo_mem[2][7] ),
	.D(n68),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][6]  (
	.SI(\fifo_mem[2][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[2][6] ),
	.D(n67),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][5]  (
	.SI(\fifo_mem[2][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[2][5] ),
	.D(n66),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][4]  (
	.SI(\fifo_mem[2][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[2][4] ),
	.D(n65),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][3]  (
	.SI(\fifo_mem[2][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[2][3] ),
	.D(n64),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][2]  (
	.SI(\fifo_mem[2][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[2][2] ),
	.D(n63),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][1]  (
	.SI(\fifo_mem[2][0] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[2][1] ),
	.D(n62),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[2][0]  (
	.SI(\fifo_mem[1][7] ),
	.SE(n122),
	.RN(wrst_n),
	.Q(\fifo_mem[2][0] ),
	.D(n61),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][7]  (
	.SI(\fifo_mem[6][6] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][7] ),
	.D(n36),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][6]  (
	.SI(\fifo_mem[6][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][6] ),
	.D(n35),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][5]  (
	.SI(\fifo_mem[6][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][5] ),
	.D(n34),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][4]  (
	.SI(\fifo_mem[6][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][4] ),
	.D(n33),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][3]  (
	.SI(\fifo_mem[6][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][3] ),
	.D(n32),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][2]  (
	.SI(\fifo_mem[6][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][2] ),
	.D(n31),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][1]  (
	.SI(\fifo_mem[6][0] ),
	.SE(n119),
	.RN(wrst_n),
	.Q(\fifo_mem[6][1] ),
	.D(n30),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[6][0]  (
	.SI(\fifo_mem[5][7] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[6][0] ),
	.D(n29),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][7]  (
	.SI(\fifo_mem[0][6] ),
	.SE(n121),
	.RN(wrst_n),
	.Q(\fifo_mem[0][7] ),
	.D(n84),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][6]  (
	.SI(\fifo_mem[0][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[0][6] ),
	.D(n83),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][5]  (
	.SI(\fifo_mem[0][4] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[0][5] ),
	.D(n82),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][4]  (
	.SI(\fifo_mem[0][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[0][4] ),
	.D(n81),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][3]  (
	.SI(\fifo_mem[0][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[0][3] ),
	.D(n80),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][2]  (
	.SI(\fifo_mem[0][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[0][2] ),
	.D(n79),
	.CK(REF_SCAN_CLK__L6_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][1]  (
	.SI(\fifo_mem[0][0] ),
	.SE(n119),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[0][1] ),
	.D(n78),
	.CK(wclk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[0][0]  (
	.SI(test_si1),
	.SE(n122),
	.RN(wrst_n),
	.Q(\fifo_mem[0][0] ),
	.D(n77),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][7]  (
	.SI(\fifo_mem[4][6] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[4][7] ),
	.D(n52),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][6]  (
	.SI(\fifo_mem[4][5] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[4][6] ),
	.D(n51),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][5]  (
	.SI(test_si2),
	.SE(n119),
	.RN(wrst_n),
	.Q(\fifo_mem[4][5] ),
	.D(n50),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][3]  (
	.SI(\fifo_mem[4][2] ),
	.SE(n121),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[4][3] ),
	.D(n48),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][2]  (
	.SI(\fifo_mem[4][1] ),
	.SE(n120),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(\fifo_mem[4][2] ),
	.D(n47),
	.CK(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][1]  (
	.SI(\fifo_mem[4][0] ),
	.SE(n119),
	.RN(wrst_n),
	.Q(\fifo_mem[4][1] ),
	.D(n46),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_mem_reg[4][0]  (
	.SI(\fifo_mem[3][7] ),
	.SE(n122),
	.RN(wrst_n),
	.Q(\fifo_mem[4][0] ),
	.D(n45),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U124 (
	.Y(n118),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U125 (
	.Y(n119),
	.A(n118), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U126 (
	.Y(n120),
	.A(n118), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U127 (
	.Y(n121),
	.A(n118), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U128 (
	.Y(n122),
	.A(n118), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U129 (
	.Y(n123),
	.A(\fifo_mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U130 (
	.Y(n124),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \fifo_mem_reg[4][4]  (
	.SI(\fifo_mem[4][3] ),
	.SE(n122),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(FE_OFN7_SO_3_),
	.D(n49),
	.CK(REF_SCAN_CLK__L6_N13), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GEN_test_1 (
	clk, 
	rst, 
	lvl_sig, 
	pulse_sig, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst;
   input lvl_sig;
   output pulse_sig;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire pls_flop;
   wire rcv_flop;

   assign test_so = rcv_flop ;

   // Module instantiations
   NOR2BX2M U3 (
	.Y(pulse_sig),
	.B(pls_flop),
	.AN(rcv_flop), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M rcv_flop_reg (
	.SI(pls_flop),
	.SE(test_se),
	.RN(rst),
	.Q(rcv_flop),
	.D(lvl_sig),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M pls_flop_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst),
	.Q(pls_flop),
	.D(rcv_flop),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	n20__Exclude_0_NET, 
	n20__L1_N0, 
	SYNC_SCAN_RST2__L1_N0, 
	UART_SCAN_CLK__L18_N0, 
	UART_SCAN_CLK__L9_N3, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input n20__Exclude_0_NET;
   input n20__L1_N0;
   input SYNC_SCAN_RST2__L1_N0;
   input UART_SCAN_CLK__L18_N0;
   input UART_SCAN_CLK__L9_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN11_n21__Exclude_0_NET;
   wire N0__L1_N0;
   wire HTIE_LTIEHI_NET;
   wire FE_UNCONNECTED_0;
   wire N0;
   wire reg_div_clk;
   wire flag;
   wire N11;
   wire N16;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire [7:0] counter;

//   assign test_so = reg_div_clk ;

   // Module instantiations
   DLY4X1M FE_PHC11_n21__Exclude_0_NET (
	.Y(FE_PHN11_n21__Exclude_0_NET),
	.A(test_si), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M N0__L1_I0 (
	.Y(N0__L1_N0),
	.A(N0), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n54),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U4 (
	.Y(N0),
	.B(n55),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U5 (
	.Y(n27),
	.B1(n57),
	.B0(n54),
	.A1(n18),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U6 (
	.Y(n18),
	.B(n19),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U7 (
	.Y(n19),
	.B0(n16),
	.A1N(N24),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n55),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n3),
	.A(SYNC_SCAN_RST2__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U10 (
	.Y(n26),
	.B1(n15),
	.B0(n14),
	.A1N(n20__Exclude_0_NET),
	.A0N(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U11 (
	.Y(n15),
	.B0(n16),
	.A1(n20__Exclude_0_NET),
	.A0(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U12 (
	.Y(n14),
	.B0(n54),
	.A2(n55),
	.A1(n56),
	.A0(N24), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U13 (
	.Y(n4),
	.B(i_div_ratio[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U14 (
	.Y(n21),
	.B(n55),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U15 (
	.Y(n22),
	.B0(n23),
	.A2(n56),
	.A1(N11),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U16 (
	.Y(n23),
	.B0(N24),
	.A1(i_div_ratio[0]),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U17 (
	.Y(n34),
	.B1(n21),
	.B0(N28),
	.A1(n20),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U18 (
	.Y(n33),
	.B1(n21),
	.B0(N29),
	.A1(n20),
	.A0(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U19 (
	.Y(n32),
	.B1(n21),
	.B0(N30),
	.A1(n20),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U20 (
	.Y(n31),
	.B1(n21),
	.B0(N31),
	.A1(n20),
	.A0(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U21 (
	.Y(n30),
	.B1(n21),
	.B0(N32),
	.A1(n20),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U22 (
	.Y(n29),
	.B1(n21),
	.B0(N33),
	.A1(n20),
	.A0(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U23 (
	.Y(n28),
	.B1(n21),
	.B0(N34),
	.A1(n20),
	.A0(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U24 (
	.Y(n35),
	.B1(n21),
	.B0(n42),
	.A1(n20),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U25 (
	.Y(n16),
	.C(flag),
	.B(i_div_ratio[0]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U26 (
	.Y(n1),
	.B0N(n4),
	.A1(i_div_ratio[2]),
	.A0(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n42),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U28 (
	.Y(n17),
	.B(n57),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n57),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U31 (
	.Y(n20),
	.B0(HTIE_LTIEHI_NET),
	.A1N(n25),
	.A0N(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U32 (
	.Y(n24),
	.C(i_div_ratio[2]),
	.B(i_div_ratio[3]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U33 (
	.Y(n25),
	.D(i_div_ratio[4]),
	.C(i_div_ratio[5]),
	.B(i_div_ratio[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n56),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U35 (
	.Y(o_div_clk),
	.S0(N0__L1_N0),
	.B(i_ref_clk),
	.A(n20__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U36 (
	.Y(N16),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U37 (
	.Y(n5),
	.B(i_div_ratio[3]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U38 (
	.Y(N18),
	.B0(n5),
	.A1N(i_div_ratio[3]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U39 (
	.Y(n6),
	.B(i_div_ratio[4]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U40 (
	.Y(N19),
	.B0(n6),
	.A1N(i_div_ratio[4]),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U41 (
	.Y(n7),
	.B(i_div_ratio[5]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U42 (
	.Y(N20),
	.B0(n7),
	.A1N(i_div_ratio[5]),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U43 (
	.Y(N21),
	.B(n7),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U44 (
	.Y(N23),
	.C(n7),
	.B(i_div_ratio[7]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U45 (
	.Y(n8),
	.B0(i_div_ratio[7]),
	.A1(n7),
	.A0(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U46 (
	.Y(N22),
	.B(n8),
	.AN(N23), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U47 (
	.Y(n41),
	.B(counter[2]),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U48 (
	.Y(n9),
	.B(N16),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U49 (
	.Y(n40),
	.B1(n1),
	.B0(n9),
	.A1(n9),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U50 (
	.Y(n10),
	.B(n42),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U51 (
	.Y(n11),
	.B1(counter[1]),
	.B0(n10),
	.A1(n1),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U52 (
	.Y(n39),
	.C(counter[7]),
	.B(N23),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U53 (
	.Y(n37),
	.B(counter[3]),
	.A(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n36),
	.B(counter[4]),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U55 (
	.Y(n13),
	.B(counter[5]),
	.A(N21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n12),
	.B(counter[6]),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U57 (
	.Y(n38),
	.D(n12),
	.C(n13),
	.B(n36),
	.A(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U58 (
	.Y(N24),
	.D(n38),
	.C(n39),
	.B(n40),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U59 (
	.Y(n43),
	.B(i_div_ratio[1]),
	.AN(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U60 (
	.Y(n47),
	.B1(n43),
	.B0(counter[1]),
	.A1N(i_div_ratio[2]),
	.A0(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U61 (
	.Y(n46),
	.B(counter[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U62 (
	.Y(n44),
	.B(counter[0]),
	.AN(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U63 (
	.Y(n45),
	.B1(n44),
	.B0(i_div_ratio[2]),
	.A1N(counter[1]),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U64 (
	.Y(n53),
	.D(n45),
	.C(n46),
	.B(n47),
	.AN(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U65 (
	.Y(n51),
	.B(counter[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U66 (
	.Y(n50),
	.B(counter[5]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U67 (
	.Y(n49),
	.B(counter[4]),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U68 (
	.Y(n48),
	.B(counter[3]),
	.A(i_div_ratio[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U69 (
	.Y(n52),
	.D(n48),
	.C(n49),
	.B(n50),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(N11),
	.B(n52),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M reg_div_clk_reg (
	.SI(n57),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(test_so),
	.D(n26),
	.CK(UART_SCAN_CLK__L9_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M flag_reg (
	.SI(counter[7]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(flag),
	.D(n27),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[7]),
	.D(n28),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(FE_PHN11_n21__Exclude_0_NET),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(n35),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(n33),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(n29),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(n30),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(n31),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(n32),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(n42),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(n34),
	.CK(UART_SCAN_CLK__L18_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_0_DW01_inc_0 r76 (
	.A({ counter[7],
		counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N34,
		N33,
		N32,
		N31,
		N30,
		N29,
		N28,
		FE_UNCONNECTED_0 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLKDIV_MUX (
	IN, 
	OUT, 
	VDD, 
	VSS);
   input [5:0] IN;
   output [7:0] OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U11 (
	.Y(OUT[0]),
	.C0(n16),
	.B0(n17),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U12 (
	.Y(OUT[1]),
	.C(IN[0]),
	.B(IN[1]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U13 (
	.Y(n6),
	.D(n14),
	.C(n15),
	.B(IN[3]),
	.AN(IN[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U14 (
	.Y(n7),
	.D(n14),
	.C(n15),
	.B(IN[4]),
	.AN(IN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(OUT[2]),
	.C(IN[0]),
	.B(IN[1]),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n15),
	.A(IN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n14),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U18 (
	.Y(OUT[3]),
	.D(IN[4]),
	.C(n19),
	.B(IN[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U19 (
	.Y(n5),
	.C(IN[2]),
	.B(n16),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n17),
	.A(IN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n16),
	.A(IN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U22 (
	.Y(n8),
	.D(n15),
	.C(IN[3]),
	.B(IN[4]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(n9),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U24 (
	.Y(n18),
	.A(IN[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U25 (
	.Y(n19),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(OUT[4]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(OUT[5]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(OUT[6]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(OUT[7]),
	.A(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_test_0 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	n21__Exclude_0_NET, 
	UART_SCAN_CLK__L18_N1, 
	UART_SCAN_CLK__L9_N2, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input n21__Exclude_0_NET;
   input UART_SCAN_CLK__L18_N1;
   input UART_SCAN_CLK__L9_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN16_n4__Exclude_0_NET;
   wire FE_PHN15_n4__Exclude_0_NET;
   wire n4__Exclude_0_NET;
   wire N0__L1_N0;
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire FE_UNCONNECTED_0;
   wire N0;
   wire reg_div_clk;
   wire flag;
   wire N11;
   wire N16;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire [7:0] counter;

//   assign test_so = reg_div_clk ;

   // Module instantiations
   DLY4X1M FE_PHC16_n4__Exclude_0_NET (
	.Y(FE_PHN15_n4__Exclude_0_NET),
	.A(FE_PHN16_n4__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC15_n4__Exclude_0_NET (
	.Y(n4__Exclude_0_NET),
	.A(FE_PHN15_n4__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M n4__Exclude_0 (
	.Y(FE_PHN16_n4__Exclude_0_NET),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M N0__L1_I0 (
	.Y(N0__L1_N0),
	.A(N0), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n55),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U4 (
	.Y(N0),
	.B(n58),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n3),
	.A(n4__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U6 (
	.Y(n76),
	.B(n75),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U7 (
	.Y(n75),
	.B0(n78),
	.A1N(N24),
	.A0(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U8 (
	.Y(n67),
	.B1(n56),
	.B0(n55),
	.A1(n76),
	.A0(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U9 (
	.Y(n5),
	.B(i_div_ratio[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U10 (
	.Y(n73),
	.B(n58),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U11 (
	.Y(n72),
	.B0(n71),
	.A2(n57),
	.A1(N11),
	.A0(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U12 (
	.Y(n71),
	.B0(N24),
	.A1(i_div_ratio[0]),
	.A0(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U13 (
	.Y(n1),
	.B0N(n5),
	.A1(i_div_ratio[2]),
	.A0(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(n77),
	.B(n56),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n57),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n58),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n4),
	.A(i_rst_n), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U18 (
	.Y(n68),
	.B1(n79),
	.B0(n80),
	.A1N(n21__Exclude_0_NET),
	.A0N(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U19 (
	.Y(n79),
	.B0(n78),
	.A1(n21__Exclude_0_NET),
	.A0(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U20 (
	.Y(n80),
	.B0(n55),
	.A2(n58),
	.A1(n57),
	.A0(N24), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U21 (
	.Y(n60),
	.B1(n73),
	.B0(N28),
	.A1(n74),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U22 (
	.Y(n61),
	.B1(n73),
	.B0(N29),
	.A1(n74),
	.A0(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U23 (
	.Y(n62),
	.B1(n73),
	.B0(N30),
	.A1(n74),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U24 (
	.Y(n63),
	.B1(n73),
	.B0(N31),
	.A1(n74),
	.A0(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n64),
	.B1(n73),
	.B0(N32),
	.A1(n74),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n65),
	.B1(n73),
	.B0(N33),
	.A1(n74),
	.A0(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n66),
	.B1(n73),
	.B0(N34),
	.A1(n74),
	.A0(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U28 (
	.Y(n59),
	.B1(n73),
	.B0(n43),
	.A1(n74),
	.A0(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U29 (
	.Y(n78),
	.C(flag),
	.B(i_div_ratio[0]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U31 (
	.Y(n74),
	.B0(HTIE_LTIEHI_NET),
	.A1N(n69),
	.A0N(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U32 (
	.Y(n69),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U33 (
	.Y(n70),
	.C(i_div_ratio[2]),
	.B(i_div_ratio[3]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n43),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U35 (
	.Y(n56),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U36 (
	.Y(o_div_clk),
	.S0(N0__L1_N0),
	.B(i_ref_clk),
	.A(test_so), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U37 (
	.Y(N16),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U38 (
	.Y(n6),
	.B(i_div_ratio[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U39 (
	.Y(N18),
	.B0(n6),
	.A1N(i_div_ratio[3]),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U40 (
	.Y(n7),
	.B(LTIE_LTIELO_NET),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U41 (
	.Y(N19),
	.B0(n7),
	.A1N(LTIE_LTIELO_NET),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U42 (
	.Y(n8),
	.B(LTIE_LTIELO_NET),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U43 (
	.Y(N20),
	.B0(n8),
	.A1N(LTIE_LTIELO_NET),
	.A0N(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U44 (
	.Y(N21),
	.B(n8),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U45 (
	.Y(N23),
	.C(n8),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U46 (
	.Y(n9),
	.B0(LTIE_LTIELO_NET),
	.A1(n8),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U47 (
	.Y(N22),
	.B(n9),
	.AN(N23), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U48 (
	.Y(n42),
	.B(counter[2]),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U49 (
	.Y(n10),
	.B(N16),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U50 (
	.Y(n41),
	.B1(n1),
	.B0(n10),
	.A1(n10),
	.A0(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U51 (
	.Y(n11),
	.B(n43),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U52 (
	.Y(n12),
	.B1(counter[1]),
	.B0(n11),
	.A1(n1),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U53 (
	.Y(n40),
	.C(counter[7]),
	.B(N23),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n38),
	.B(counter[3]),
	.A(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U55 (
	.Y(n37),
	.B(counter[4]),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n36),
	.B(counter[5]),
	.A(N21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n13),
	.B(counter[6]),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U58 (
	.Y(n39),
	.D(n13),
	.C(n36),
	.B(n37),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U59 (
	.Y(N24),
	.D(n39),
	.C(n40),
	.B(n41),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U60 (
	.Y(n44),
	.B(i_div_ratio[1]),
	.AN(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U61 (
	.Y(n48),
	.B1(n44),
	.B0(counter[1]),
	.A1N(i_div_ratio[2]),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U62 (
	.Y(n47),
	.B(counter[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U63 (
	.Y(n45),
	.B(counter[0]),
	.AN(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U64 (
	.Y(n46),
	.B1(n45),
	.B0(i_div_ratio[2]),
	.A1N(counter[1]),
	.A0(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U65 (
	.Y(n54),
	.D(n46),
	.C(n47),
	.B(n48),
	.AN(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U66 (
	.Y(n52),
	.B(counter[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U67 (
	.Y(n51),
	.B(counter[5]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U68 (
	.Y(n50),
	.B(counter[4]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U69 (
	.Y(n49),
	.B(counter[3]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U70 (
	.Y(n53),
	.D(n49),
	.C(n50),
	.B(n51),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(N11),
	.B(n53),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M reg_div_clk_reg (
	.SI(n56),
	.SE(test_se),
	.RN(n3),
	.Q(test_so),
	.D(n68),
	.CK(UART_SCAN_CLK__L9_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M flag_reg (
	.SI(counter[7]),
	.SE(test_se),
	.RN(n3),
	.Q(flag),
	.D(n67),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(n3),
	.Q(counter[7]),
	.D(n66),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(n3),
	.Q(counter[0]),
	.D(n59),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(n3),
	.Q(counter[2]),
	.D(n61),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(n3),
	.Q(counter[6]),
	.D(n65),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(n3),
	.Q(counter[5]),
	.D(n64),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(n3),
	.Q(counter[4]),
	.D(n63),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(n3),
	.Q(counter[3]),
	.D(n62),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(n43),
	.SE(test_se),
	.RN(n3),
	.Q(counter[1]),
	.D(n60),
	.CK(UART_SCAN_CLK__L18_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_1_DW01_inc_0 r76 (
	.A({ counter[7],
		counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N34,
		N33,
		N32,
		N31,
		N30,
		N29,
		N28,
		FE_UNCONNECTED_0 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ClkDiv_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_DATA_WIDTH8_test_1 (
	RST, 
	TX_CLK, 
	RX_CLK, 
	RX_IN_S, 
	RX_OUT_P, 
	RX_OUT_V, 
	TX_IN_P, 
	TX_IN_V, 
	TX_OUT_S, 
	TX_OUT_V, 
	Prescale, 
	parity_enable, 
	parity_type, 
	parity_error, 
	framing_error, 
	test_si, 
	test_se, 
	TX_SCAN_CLK__L4_N1, 
	RX_SCAN_CLK__L4_N1, 
	VDD, 
	VSS);
   input RST;
   input TX_CLK;
   input RX_CLK;
   input RX_IN_S;
   output [7:0] RX_OUT_P;
   output RX_OUT_V;
   input [7:0] TX_IN_P;
   input TX_IN_V;
   output TX_OUT_S;
   output TX_OUT_V;
   input [5:0] Prescale;
   input parity_enable;
   input parity_type;
   output parity_error;
   output framing_error;
   input test_si;
   input test_se;
   input TX_SCAN_CLK__L4_N1;
   input RX_SCAN_CLK__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;

   // Module instantiations
   UART_TX_DATA_WIDTH8_test_1 U0_UART_TX (
	.CLK(TX_CLK),
	.RST(RST),
	.P_DATA({ TX_IN_P[7],
		TX_IN_P[6],
		TX_IN_P[5],
		TX_IN_P[4],
		TX_IN_P[3],
		TX_IN_P[2],
		TX_IN_P[1],
		TX_IN_P[0] }),
	.Data_Valid(TX_IN_V),
	.parity_enable(parity_enable),
	.parity_type(parity_type),
	.TX_OUT(TX_OUT_S),
	.busy(TX_OUT_V),
	.test_si(n3),
	.test_se(test_se),
	.TX_SCAN_CLK__L4_N1(TX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_RX_test_1 U0_UART_RX (
	.CLK(RX_CLK),
	.RST(RST),
	.RX_IN(RX_IN_S),
	.parity_enable(parity_enable),
	.parity_type(parity_type),
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.P_DATA({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.data_valid(RX_OUT_V),
	.parity_error(parity_error),
	.framing_error(framing_error),
	.test_si(test_si),
	.test_so(n3),
	.test_se(test_se),
	.RX_SCAN_CLK__L4_N1(RX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_TX_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	P_DATA, 
	Data_Valid, 
	parity_enable, 
	parity_type, 
	TX_OUT, 
	busy, 
	test_si, 
	test_se, 
	TX_SCAN_CLK__L4_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] P_DATA;
   input Data_Valid;
   input parity_enable;
   input parity_type;
   output TX_OUT;
   output busy;
   input test_si;
   input test_se;
   input TX_SCAN_CLK__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire seriz_done;
   wire seriz_en;
   wire ser_data;
   wire parity;
   wire n3;
   wire n4;
   wire [1:0] mux_sel;

   // Module instantiations
   uart_tx_fsm_test_1 U0_fsm (
	.CLK(TX_SCAN_CLK__L4_N1),
	.RST(RST),
	.Data_Valid(Data_Valid),
	.ser_done(seriz_done),
	.parity_enable(parity_enable),
	.Ser_enable(seriz_en),
	.mux_sel({ mux_sel[1],
		mux_sel[0] }),
	.busy(busy),
	.test_si(n4),
	.test_so(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   Serializer_WIDTH8_test_1 U0_Serializer (
	.CLK(TX_SCAN_CLK__L4_N1),
	.RST(RST),
	.DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.Enable(seriz_en),
	.Busy(busy),
	.Data_Valid(Data_Valid),
	.ser_out(ser_data),
	.ser_done(seriz_done),
	.test_si(test_si),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_test_1 U0_mux (
	.CLK(CLK),
	.RST(RST),
	.IN_0(1'b0),
	.IN_1(ser_data),
	.IN_2(parity),
	.IN_3(1'b1),
	.SEL({ mux_sel[1],
		mux_sel[0] }),
	.OUT(TX_OUT),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_calc_WIDTH8_test_1 U0_parity_calc (
	.CLK(CLK),
	.RST(RST),
	.parity_enable(parity_enable),
	.parity_type(parity_type),
	.Busy(busy),
	.DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.Data_Valid(Data_Valid),
	.parity(parity),
	.test_si(n3),
	.test_se(test_se),
	.TX_SCAN_CLK__L4_N1(TX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module uart_tx_fsm_test_1 (
	CLK, 
	RST, 
	Data_Valid, 
	ser_done, 
	parity_enable, 
	Ser_enable, 
	mux_sel, 
	busy, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input Data_Valid;
   input ser_done;
   input parity_enable;
   output Ser_enable;
   output [1:0] mux_sel;
   output busy;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire busy_c;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n1;
   wire n2;
   wire n3;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   // Module instantiations
   INVX2M U3 (
	.Y(n1),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U4 (
	.Y(Ser_enable),
	.C(current_state[2]),
	.B(ser_done),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U5 (
	.Y(n9),
	.B0(n8),
	.A1(n2),
	.A0(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U6 (
	.Y(n8),
	.B(n2),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n5),
	.B(current_state[0]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n2),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U9 (
	.Y(mux_sel[0]),
	.B1(n9),
	.B0(current_state[2]),
	.A1N(current_state[2]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U10 (
	.Y(mux_sel[1]),
	.B0(n8),
	.A1(current_state[0]),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U11 (
	.Y(next_state[2]),
	.C(n4),
	.B(current_state[2]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U12 (
	.Y(n4),
	.B0(n2),
	.A1N(parity_enable),
	.A0(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U13 (
	.Y(busy_c),
	.B0(n8),
	.A1(n2),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U14 (
	.Y(next_state[1]),
	.B0(current_state[2]),
	.A1(n5),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U15 (
	.Y(next_state[0]),
	.B0(current_state[2]),
	.A1(n7),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U16 (
	.Y(n6),
	.B(current_state[0]),
	.AN(ser_done), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U17 (
	.Y(n7),
	.B0(n3),
	.A1(current_state[0]),
	.A0(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n3),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M busy_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(busy),
	.D(busy_c),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n3),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(busy),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Serializer_WIDTH8_test_1 (
	CLK, 
	RST, 
	DATA, 
	Enable, 
	Busy, 
	Data_Valid, 
	ser_out, 
	ser_done, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] DATA;
   input Enable;
   input Busy;
   input Data_Valid;
   output ser_out;
   output ser_done;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N23;
   wire N24;
   wire N25;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n2;
   wire n3;
   wire n25;
   wire n28;
   wire n29;
   wire [7:1] DATA_V;
   wire [2:0] ser_count;

   assign test_so = n25 ;

   // Module instantiations
   NOR2X2M U3 (
	.Y(n6),
	.B(n7),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U4 (
	.Y(n4),
	.B(n6),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n2),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U6 (
	.Y(N25),
	.B1(n25),
	.B0(n15),
	.A2(n2),
	.A1(n3),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n14),
	.B(n25),
	.A(ser_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U8 (
	.Y(n15),
	.B0(N23),
	.A1(n3),
	.A0(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n25),
	.A(ser_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U11 (
	.Y(n7),
	.B(Busy),
	.AN(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U12 (
	.Y(n17),
	.B0(n5),
	.A1N(n4),
	.A0N(ser_out), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U13 (
	.Y(n5),
	.B1(n7),
	.B0(DATA[0]),
	.A1(n6),
	.A0(DATA_V[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U14 (
	.Y(n24),
	.B0(n13),
	.A1N(n4),
	.A0N(DATA_V[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U15 (
	.Y(n13),
	.B1(n7),
	.B0(DATA[1]),
	.A1(n6),
	.A0(DATA_V[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U16 (
	.Y(n23),
	.B0(n12),
	.A1N(DATA_V[2]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U17 (
	.Y(n12),
	.B1(n7),
	.B0(DATA[2]),
	.A1(n6),
	.A0(DATA_V[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U18 (
	.Y(n22),
	.B0(n11),
	.A1N(DATA_V[3]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U19 (
	.Y(n11),
	.B1(n7),
	.B0(DATA[3]),
	.A1(n6),
	.A0(DATA_V[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U20 (
	.Y(n21),
	.B0(n10),
	.A1N(DATA_V[4]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U21 (
	.Y(n10),
	.B1(n7),
	.B0(DATA[4]),
	.A1(n6),
	.A0(DATA_V[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U22 (
	.Y(n20),
	.B0(n9),
	.A1N(DATA_V[5]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U23 (
	.Y(n9),
	.B1(n7),
	.B0(DATA[5]),
	.A1(n6),
	.A0(DATA_V[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U24 (
	.Y(n19),
	.B0(n8),
	.A1N(DATA_V[6]),
	.A0N(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U25 (
	.Y(n8),
	.B1(n7),
	.B0(DATA[6]),
	.A1(n6),
	.A0(DATA_V[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n18),
	.B1(n7),
	.B0(DATA[7]),
	.A1(DATA_V[7]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U27 (
	.Y(ser_done),
	.C(ser_count[1]),
	.B(ser_count[2]),
	.A(ser_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U28 (
	.Y(N23),
	.B(ser_count[0]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(N24),
	.B(n2),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n16),
	.B(n3),
	.A(ser_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n3),
	.A(ser_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[0]  (
	.SI(test_si),
	.SE(n29),
	.RN(RST),
	.Q(ser_out),
	.D(n17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[6]  (
	.SI(DATA_V[5]),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[6]),
	.D(n19),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[5]  (
	.SI(DATA_V[4]),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[5]),
	.D(n20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[4]  (
	.SI(DATA_V[3]),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[4]),
	.D(n21),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[3]  (
	.SI(DATA_V[2]),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[3]),
	.D(n22),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[2]  (
	.SI(DATA_V[1]),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[2]),
	.D(n23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[1]  (
	.SI(ser_out),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[1]),
	.D(n24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[7]  (
	.SI(DATA_V[6]),
	.SE(n29),
	.RN(RST),
	.Q(DATA_V[7]),
	.D(n18),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ser_count_reg[2]  (
	.SI(n3),
	.SE(n29),
	.RN(RST),
	.Q(ser_count[2]),
	.D(N25),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ser_count_reg[1]  (
	.SI(ser_count[0]),
	.SE(n29),
	.RN(RST),
	.Q(ser_count[1]),
	.D(N24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ser_count_reg[0]  (
	.SI(DATA_V[7]),
	.SE(n29),
	.RN(RST),
	.Q(ser_count[0]),
	.D(N23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U32 (
	.Y(n28),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U33 (
	.Y(n29),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_test_1 (
	CLK, 
	RST, 
	IN_0, 
	IN_1, 
	IN_2, 
	IN_3, 
	SEL, 
	OUT, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input IN_0;
   input IN_1;
   input IN_2;
   input IN_3;
   input [1:0] SEL;
   output OUT;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire mux_out;
   wire n2;
   wire n3;
   wire n1;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n1),
	.A(SEL[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U4 (
	.Y(mux_out),
	.B1(n3),
	.B0(SEL[1]),
	.A1N(SEL[1]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U5 (
	.Y(n3),
	.B1(IN_1),
	.B0(SEL[0]),
	.A1(n1),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U6 (
	.Y(n2),
	.B1(SEL[0]),
	.B0(HTIE_LTIEHI_NET),
	.A1(n1),
	.A0(IN_2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M OUT_reg (
	.SI(IN_2),
	.SE(test_se),
	.RN(RST),
	.Q(OUT),
	.D(mux_out),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_calc_WIDTH8_test_1 (
	CLK, 
	RST, 
	parity_enable, 
	parity_type, 
	Busy, 
	DATA, 
	Data_Valid, 
	parity, 
	test_si, 
	test_se, 
	TX_SCAN_CLK__L4_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input parity_enable;
   input parity_type;
   input Busy;
   input [7:0] DATA;
   input Data_Valid;
   output parity;
   input test_si;
   input test_se;
   input TX_SCAN_CLK__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n2;
   wire [7:0] DATA_V;

   // Module instantiations
   NOR2BX2M U2 (
	.Y(n7),
	.B(Busy),
	.AN(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U3 (
	.Y(n9),
	.B1(n7),
	.B0(DATA[0]),
	.A1N(n7),
	.A0(DATA_V[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U4 (
	.Y(n10),
	.B1(n7),
	.B0(DATA[1]),
	.A1N(n7),
	.A0(DATA_V[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U5 (
	.Y(n11),
	.B1(n7),
	.B0(DATA[2]),
	.A1N(n7),
	.A0(DATA_V[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U6 (
	.Y(n12),
	.B1(n7),
	.B0(DATA[3]),
	.A1N(n7),
	.A0(DATA_V[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U7 (
	.Y(n13),
	.B1(n7),
	.B0(DATA[4]),
	.A1N(n7),
	.A0(DATA_V[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U8 (
	.Y(n14),
	.B1(n7),
	.B0(DATA[5]),
	.A1N(n7),
	.A0(DATA_V[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U9 (
	.Y(n15),
	.B1(n7),
	.B0(DATA[6]),
	.A1N(n7),
	.A0(DATA_V[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U10 (
	.Y(n16),
	.B1(n7),
	.B0(DATA[7]),
	.A1N(n7),
	.A0(DATA_V[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U11 (
	.Y(n5),
	.B(DATA_V[3]),
	.A(DATA_V[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(n8),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(parity), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n2),
	.A(parity_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U14 (
	.Y(n1),
	.C(n4),
	.B(parity_type),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U15 (
	.Y(n4),
	.C(n5),
	.B(DATA_V[0]),
	.A(DATA_V[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U16 (
	.Y(n3),
	.C(n6),
	.B(DATA_V[4]),
	.A(DATA_V[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(n6),
	.B(DATA_V[6]),
	.A(DATA_V[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M parity_reg (
	.SI(DATA_V[7]),
	.SE(test_se),
	.RN(RST),
	.Q(parity),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[5]  (
	.SI(DATA_V[4]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[5]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[1]  (
	.SI(DATA_V[0]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[1]),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[4]  (
	.SI(DATA_V[3]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[4]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[0]),
	.D(n9),
	.CK(TX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[2]  (
	.SI(DATA_V[1]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[2]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[3]  (
	.SI(DATA_V[2]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[3]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[6]  (
	.SI(DATA_V[5]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[6]),
	.D(n15),
	.CK(TX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \DATA_V_reg[7]  (
	.SI(DATA_V[6]),
	.SE(test_se),
	.RN(RST),
	.Q(DATA_V[7]),
	.D(n16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_RX_test_1 (
	CLK, 
	RST, 
	RX_IN, 
	parity_enable, 
	parity_type, 
	Prescale, 
	P_DATA, 
	data_valid, 
	parity_error, 
	framing_error, 
	test_si, 
	test_so, 
	test_se, 
	RX_SCAN_CLK__L4_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input RX_IN;
   input parity_enable;
   input parity_type;
   input [5:0] Prescale;
   output [7:0] P_DATA;
   output data_valid;
   output parity_error;
   output framing_error;
   input test_si;
   output test_so;
   input test_se;
   input RX_SCAN_CLK__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n15;
   wire n16;
   wire strt_glitch;
   wire strt_chk_en;
   wire edge_bit_en;
   wire deser_en;
   wire par_chk_en;
   wire stp_chk_en;
   wire dat_samp_en;
   wire sampled_bit;
   wire n4;
   wire n13;
   wire n14;
   wire [3:0] bit_count;
   wire [5:0] edge_count;

   // Module instantiations
   INVXLM U9 (
	.Y(n13),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U10 (
	.Y(n14),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   uart_rx_fsm_DATA_WIDTH8_test_1 U0_uart_fsm (
	.CLK(CLK),
	.RST(RST),
	.S_DATA(RX_IN),
	.Prescale({ n14,
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.parity_enable(parity_enable),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.par_err(n15),
	.stp_err(n16),
	.strt_glitch(strt_glitch),
	.strt_chk_en(strt_chk_en),
	.edge_bit_en(edge_bit_en),
	.deser_en(deser_en),
	.par_chk_en(par_chk_en),
	.stp_chk_en(stp_chk_en),
	.dat_samp_en(dat_samp_en),
	.data_valid(data_valid),
	.test_so(test_so),
	.test_se(test_se),
	.RX_SCAN_CLK__L4_N1(RX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   edge_bit_counter_test_1 U0_edge_bit_counter (
	.CLK(RX_SCAN_CLK__L4_N1),
	.RST(RST),
	.Enable(edge_bit_en),
	.Prescale({ n14,
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.bit_count({ bit_count[3],
		bit_count[2],
		bit_count[1],
		bit_count[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.test_si(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   data_sampling_test_1 U0_data_sampling (
	.CLK(CLK),
	.RST(RST),
	.S_DATA(RX_IN),
	.Prescale({ n14,
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.Enable(dat_samp_en),
	.sampled_bit(sampled_bit),
	.test_si(test_si),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_DATA_WIDTH8_test_1 U0_deserializer (
	.CLK(CLK),
	.RST(RST),
	.sampled_bit(sampled_bit),
	.Enable(deser_en),
	.edge_count({ edge_count[5],
		edge_count[4],
		edge_count[3],
		edge_count[2],
		edge_count[1],
		edge_count[0] }),
	.Prescale({ n14,
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   strt_chk_test_1 U0_strt_chk (
	.CLK(RX_SCAN_CLK__L4_N1),
	.RST(RST),
	.sampled_bit(sampled_bit),
	.Enable(strt_chk_en),
	.strt_glitch(strt_glitch),
	.test_si(n16),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   par_chk_DATA_WIDTH8_test_1 U0_par_chk (
	.CLK(CLK),
	.RST(RST),
	.parity_type(parity_type),
	.sampled_bit(sampled_bit),
	.Enable(par_chk_en),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.par_err(n15),
	.test_si(edge_count[5]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   stp_chk_test_1 U0_stp_chk (
	.CLK(CLK),
	.RST(RST),
	.sampled_bit(sampled_bit),
	.Enable(stp_chk_en),
	.stp_err(n16),
	.test_si(n15),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M U3 (
	.Y(parity_error),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M U6 (
	.Y(framing_error),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module uart_rx_fsm_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	S_DATA, 
	Prescale, 
	parity_enable, 
	bit_count, 
	edge_count, 
	par_err, 
	stp_err, 
	strt_glitch, 
	strt_chk_en, 
	edge_bit_en, 
	deser_en, 
	par_chk_en, 
	stp_chk_en, 
	dat_samp_en, 
	data_valid, 
	test_so, 
	test_se, 
	RX_SCAN_CLK__L4_N1, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input S_DATA;
   input [5:0] Prescale;
   input parity_enable;
   input [3:0] bit_count;
   input [5:0] edge_count;
   input par_err;
   input stp_err;
   input strt_glitch;
   output strt_chk_en;
   output edge_bit_en;
   output deser_en;
   output par_chk_en;
   output stp_chk_en;
   output dat_samp_en;
   output data_valid;
   output test_so;
   input test_se;
   input RX_SCAN_CLK__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \sub_41/carry[5] ;
   wire \sub_41/carry[4] ;
   wire \sub_41/carry[3] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire [5:0] check_edge;
   wire [5:0] error_check_edge;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign error_check_edge[0] = Prescale[0] ;
   assign test_so = n22 ;

   // Module instantiations
   NOR3XLM U3 (
	.Y(data_valid),
	.C(par_err),
	.B(stp_err),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U4 (
	.Y(n1),
	.B(error_check_edge[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n5),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(n34),
	.B(edge_count[1]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U7 (
	.Y(error_check_edge[5]),
	.B(\sub_41/carry[5] ),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U8 (
	.Y(\sub_41/carry[5] ),
	.B(\sub_41/carry[4] ),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U9 (
	.Y(error_check_edge[4]),
	.B(Prescale[4]),
	.A(\sub_41/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U10 (
	.Y(\sub_41/carry[4] ),
	.B(\sub_41/carry[3] ),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U11 (
	.Y(error_check_edge[3]),
	.B(Prescale[3]),
	.A(\sub_41/carry[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U12 (
	.Y(\sub_41/carry[3] ),
	.B(Prescale[1]),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U13 (
	.Y(error_check_edge[2]),
	.B(Prescale[2]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U14 (
	.Y(check_edge[0]),
	.A(error_check_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U15 (
	.Y(check_edge[1]),
	.B0(n1),
	.A1N(Prescale[1]),
	.A0N(error_check_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n2),
	.B(Prescale[2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U17 (
	.Y(check_edge[2]),
	.B0(n2),
	.A1(Prescale[2]),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U18 (
	.Y(n3),
	.B(n5),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(check_edge[3]),
	.B0(n3),
	.A1(n5),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U20 (
	.Y(check_edge[4]),
	.B(n3),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U21 (
	.Y(n4),
	.B(n3),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(check_edge[5]),
	.B(n4),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U23 (
	.Y(strt_chk_en),
	.B(n6),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(par_chk_en),
	.B(n7),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U25 (
	.Y(next_state[2]),
	.B0(n10),
	.A2(n9),
	.A1(parity_enable),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U26 (
	.Y(n10),
	.B0(stp_chk_en),
	.A2(n13),
	.A1(n12),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U27 (
	.Y(n13),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U28 (
	.Y(n15),
	.A(bit_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U29 (
	.Y(n12),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U30 (
	.Y(next_state[1]),
	.B0(n7),
	.A1(n16),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U31 (
	.Y(n16),
	.B0(current_state[1]),
	.A2(n17),
	.A1(n11),
	.A0(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U32 (
	.Y(n17),
	.C(bit_count[3]),
	.B(strt_glitch),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U33 (
	.Y(next_state[0]),
	.C0(n20),
	.B1(n8),
	.B0(n19),
	.A1(n18),
	.A0(S_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U34 (
	.Y(n20),
	.B0(n24),
	.A2(n23),
	.A1(n22),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U35 (
	.Y(n24),
	.D(n28),
	.C(n27),
	.B(n26),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(n28),
	.B(edge_count[5]),
	.A(error_check_edge[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n27),
	.B(edge_count[4]),
	.A(error_check_edge[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX1M U38 (
	.Y(n26),
	.C(stp_chk_en),
	.B(bit_count[3]),
	.AN(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U39 (
	.Y(stp_chk_en),
	.B(n7),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U40 (
	.Y(n25),
	.D(n32),
	.C(n31),
	.B(n30),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U41 (
	.Y(n32),
	.B(error_check_edge[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U42 (
	.Y(n31),
	.B(n34),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n33),
	.B(edge_count[0]),
	.A(error_check_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U44 (
	.Y(n30),
	.B(error_check_edge[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U45 (
	.Y(n29),
	.S0(parity_enable),
	.B(n36),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U46 (
	.Y(n36),
	.B(n14),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U47 (
	.Y(n35),
	.B(n14),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U48 (
	.Y(n23),
	.S0(current_state[0]),
	.B(n37),
	.A(S_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U49 (
	.Y(n37),
	.D(n38),
	.C(bit_count[0]),
	.B(bit_count[3]),
	.AN(strt_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U50 (
	.Y(n19),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U51 (
	.Y(n9),
	.C(bit_count[3]),
	.B(n14),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U52 (
	.Y(n14),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U53 (
	.Y(n11),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U54 (
	.Y(n38),
	.B(n40),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U55 (
	.Y(n40),
	.D(n42),
	.C(n41),
	.B(bit_count[1]),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n42),
	.B(check_edge[0]),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n41),
	.B(check_edge[4]),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U58 (
	.Y(n39),
	.D(n46),
	.C(n45),
	.B(n44),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n46),
	.B(check_edge[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U60 (
	.Y(n45),
	.B(check_edge[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U61 (
	.Y(n44),
	.B(check_edge[5]),
	.A(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U62 (
	.Y(n43),
	.B(check_edge[1]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U63 (
	.Y(edge_bit_en),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U64 (
	.Y(n7),
	.B(n47),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U65 (
	.Y(deser_en),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U66 (
	.Y(n8),
	.C(current_state[0]),
	.B(n22),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U67 (
	.Y(n22),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U68 (
	.Y(n18),
	.C(current_state[0]),
	.B(current_state[1]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U69 (
	.Y(dat_samp_en),
	.B(n6),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U70 (
	.Y(n6),
	.B0(current_state[2]),
	.A1(S_DATA),
	.A0(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U71 (
	.Y(n47),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U72 (
	.Y(n21),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n21),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(strt_glitch),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(RX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(RX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module edge_bit_counter_test_1 (
	CLK, 
	RST, 
	Enable, 
	Prescale, 
	bit_count, 
	edge_count, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input Enable;
   input [5:0] Prescale;
   output [3:0] bit_count;
   output [5:0] edge_count;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire n4;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire \add_31/carry[5] ;
   wire \add_31/carry[4] ;
   wire \add_31/carry[3] ;
   wire \add_31/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n36;
   wire n37;

   // Module instantiations
   INVX2M U3 (
	.Y(n29),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n33),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(n13),
	.B(N31),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U6 (
	.Y(n16),
	.B0(n13),
	.A1(Enable),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U7 (
	.Y(N20),
	.B(n29),
	.AN(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U8 (
	.Y(N21),
	.B(n29),
	.AN(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U9 (
	.Y(N22),
	.B(n29),
	.AN(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U10 (
	.Y(N23),
	.B(n29),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U11 (
	.Y(n20),
	.B1(n29),
	.B0(n30),
	.A2(n13),
	.A1(bit_count[0]),
	.A0(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U12 (
	.Y(n18),
	.B1(n32),
	.B0(n15),
	.A2(n31),
	.A1(bit_count[2]),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U13 (
	.Y(n15),
	.B0N(n16),
	.A1(n31),
	.A0(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U14 (
	.Y(n17),
	.B1(n4),
	.B0(n11),
	.A2(n33),
	.A1(n10),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U16 (
	.Y(n9),
	.C(bit_count[2]),
	.B(n4),
	.A(N31), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X2M U17 (
	.Y(n12),
	.B0(n33),
	.A1N(n32),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U18 (
	.Y(n14),
	.C(Enable),
	.B(n29),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U19 (
	.Y(n19),
	.B1(n14),
	.B0(bit_count[1]),
	.A1(n31),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U20 (
	.Y(n2),
	.B(Prescale[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(N24),
	.B(n29),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U22 (
	.Y(n1),
	.B(edge_count[5]),
	.A(\add_31/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(N19),
	.B(n29),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n7),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(n10),
	.B(bit_count[0]),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n30),
	.A(bit_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n31),
	.A(bit_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U28 (
	.S(N8),
	.CO(\add_31/carry[2] ),
	.B(edge_count[0]),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U29 (
	.S(N9),
	.CO(\add_31/carry[3] ),
	.B(\add_31/carry[2] ),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U30 (
	.S(N10),
	.CO(\add_31/carry[4] ),
	.B(\add_31/carry[3] ),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n32),
	.A(bit_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U32 (
	.S(N11),
	.CO(\add_31/carry[5] ),
	.B(\add_31/carry[4] ),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U33 (
	.Y(N25),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U34 (
	.Y(N26),
	.B0(n2),
	.A1N(Prescale[1]),
	.A0N(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U35 (
	.Y(n3),
	.B(Prescale[2]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U36 (
	.Y(N27),
	.B0(n3),
	.A1(Prescale[2]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U37 (
	.Y(n5),
	.B(n7),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U38 (
	.Y(N28),
	.B0(n5),
	.A1(n7),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U39 (
	.Y(N29),
	.B(n5),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U40 (
	.Y(n6),
	.B(n5),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(N30),
	.B(n6),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U42 (
	.Y(n8),
	.B(N25),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U43 (
	.Y(n24),
	.B1(n8),
	.B0(edge_count[1]),
	.A1N(N26),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U44 (
	.Y(n21),
	.B(edge_count[0]),
	.AN(N25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U45 (
	.Y(n23),
	.B1(n21),
	.B0(N26),
	.A1N(edge_count[1]),
	.A0(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U46 (
	.Y(n22),
	.B(edge_count[5]),
	.A(N30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U47 (
	.Y(n28),
	.C(n22),
	.B(n23),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n27),
	.B(edge_count[4]),
	.A(N29), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n26),
	.B(edge_count[2]),
	.A(N27), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n25),
	.B(edge_count[3]),
	.A(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U51 (
	.Y(N31),
	.D(n25),
	.C(n26),
	.B(n27),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \bit_count_reg[3]  (
	.SI(n32),
	.SE(n37),
	.RN(RST),
	.QN(n4),
	.Q(bit_count[3]),
	.D(n17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[2]  (
	.SI(n31),
	.SE(n37),
	.RN(RST),
	.Q(bit_count[2]),
	.D(n18),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[1]  (
	.SI(n30),
	.SE(n37),
	.RN(RST),
	.Q(bit_count[1]),
	.D(n19),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_count_reg[0]  (
	.SI(test_si),
	.SE(n37),
	.RN(RST),
	.Q(bit_count[0]),
	.D(n20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[5]  (
	.SI(edge_count[4]),
	.SE(n37),
	.RN(RST),
	.Q(edge_count[5]),
	.D(N24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[4]  (
	.SI(edge_count[3]),
	.SE(n37),
	.RN(RST),
	.Q(edge_count[4]),
	.D(N23),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[3]  (
	.SI(edge_count[2]),
	.SE(n37),
	.RN(RST),
	.Q(edge_count[3]),
	.D(N22),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[2]  (
	.SI(edge_count[1]),
	.SE(n37),
	.RN(RST),
	.Q(edge_count[2]),
	.D(N21),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[1]  (
	.SI(edge_count[0]),
	.SE(n37),
	.RN(RST),
	.Q(edge_count[1]),
	.D(N20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_count_reg[0]  (
	.SI(n4),
	.SE(n37),
	.RN(RST),
	.Q(edge_count[0]),
	.D(N19),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U52 (
	.Y(n36),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U53 (
	.Y(n37),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampling_test_1 (
	CLK, 
	RST, 
	S_DATA, 
	Prescale, 
	edge_count, 
	Enable, 
	sampled_bit, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input S_DATA;
   input [5:0] Prescale;
   input [5:0] edge_count;
   input Enable;
   output sampled_bit;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N58;
   wire n19;
   wire n20;
   wire n21;
   wire \add_21/carry[4] ;
   wire \add_21/carry[3] ;
   wire \add_21/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire [4:0] half_edges;
   wire [4:0] half_edges_p1;
   wire [4:0] half_edges_n1;
   wire [2:0] Samples;

   // Module instantiations
   INVX2M U3 (
	.Y(n8),
	.A(half_edges[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U4 (
	.S(half_edges_p1[2]),
	.CO(\add_21/carry[3] ),
	.B(\add_21/carry[2] ),
	.A(half_edges[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U5 (
	.S(half_edges_p1[1]),
	.CO(\add_21/carry[2] ),
	.B(half_edges[0]),
	.A(half_edges[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U6 (
	.S(half_edges_p1[3]),
	.CO(\add_21/carry[4] ),
	.B(\add_21/carry[3] ),
	.A(half_edges[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n4),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U8 (
	.Y(half_edges[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U9 (
	.Y(n1),
	.B(Prescale[1]),
	.A(Prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U10 (
	.Y(half_edges[1]),
	.B0(n1),
	.A1(Prescale[2]),
	.A0(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U11 (
	.Y(n2),
	.B(n4),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U12 (
	.Y(half_edges[2]),
	.B0(n2),
	.A1(n4),
	.A0(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U13 (
	.Y(half_edges[3]),
	.B(n2),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U14 (
	.Y(n3),
	.B(n2),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(half_edges[4]),
	.B(n3),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(half_edges_p1[4]),
	.B(half_edges[4]),
	.A(\add_21/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U17 (
	.Y(n5),
	.B(half_edges[0]),
	.A(half_edges[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U18 (
	.Y(half_edges_n1[1]),
	.B0(n5),
	.A1(half_edges[1]),
	.A0(half_edges[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U19 (
	.Y(n6),
	.B(n8),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U20 (
	.Y(half_edges_n1[2]),
	.B0(n6),
	.A1(n8),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U21 (
	.Y(half_edges_n1[3]),
	.B(n6),
	.A(half_edges[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U22 (
	.Y(n7),
	.B(n6),
	.A(half_edges[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(half_edges_n1[4]),
	.B(n7),
	.A(half_edges[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U24 (
	.Y(n21),
	.S0(n11),
	.B(n10),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U25 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U26 (
	.Y(n13),
	.D(n17),
	.C(n16),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(n17),
	.B(half_edges_p1[1]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U28 (
	.Y(n16),
	.B(half_edges_p1[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U29 (
	.Y(n15),
	.B(half_edges_p1[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n14),
	.B(half_edges_p1[4]),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U31 (
	.Y(n12),
	.D(n25),
	.C(n24),
	.B(n23),
	.AN(edge_count[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U32 (
	.Y(n23),
	.B(Prescale[1]),
	.A(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U33 (
	.Y(n9),
	.B(Enable),
	.A(Samples[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U34 (
	.Y(n20),
	.S0(n24),
	.B(n26),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U35 (
	.Y(n24),
	.D(n30),
	.C(n29),
	.B(n28),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U36 (
	.Y(n30),
	.D(n32),
	.C(n31),
	.B(edge_count[5]),
	.AN(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n32),
	.B(edge_count[1]),
	.A(half_edges[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n31),
	.B(edge_count[0]),
	.A(half_edges[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U39 (
	.Y(n29),
	.B(half_edges[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n28),
	.B(half_edges[4]),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U41 (
	.Y(n22),
	.A(edge_count[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U42 (
	.Y(n27),
	.B(half_edges[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U43 (
	.Y(n26),
	.B(Enable),
	.A(Samples[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U44 (
	.Y(n19),
	.S0(n25),
	.B(n33),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U45 (
	.Y(n25),
	.D(n37),
	.C(n36),
	.B(n35),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U46 (
	.Y(n37),
	.C(n39),
	.B(edge_count[5]),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U47 (
	.Y(n39),
	.B(edge_count[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n38),
	.B(edge_count[4]),
	.A(half_edges_n1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U49 (
	.Y(n36),
	.B(half_edges_n1[2]),
	.A(edge_count[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U50 (
	.Y(n35),
	.B(half_edges_n1[3]),
	.A(edge_count[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n34),
	.B(half_edges_n1[1]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U52 (
	.Y(n18),
	.A(edge_count[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U53 (
	.Y(n33),
	.B(Enable),
	.A(Samples[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U54 (
	.Y(n10),
	.B(Enable),
	.A(S_DATA), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX1M U55 (
	.Y(N58),
	.B0N(Enable),
	.A1(n41),
	.A0(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U56 (
	.Y(n41),
	.B0(Samples[2]),
	.A1(Samples[1]),
	.A0(Samples[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U57 (
	.Y(n40),
	.B(Samples[1]),
	.A(Samples[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Samples_reg[2]  (
	.SI(Samples[1]),
	.SE(test_se),
	.RN(RST),
	.Q(Samples[2]),
	.D(n21),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Samples_reg[1]  (
	.SI(Samples[0]),
	.SE(test_se),
	.RN(RST),
	.Q(Samples[1]),
	.D(n20),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Samples_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(Samples[0]),
	.D(n19),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sampled_bit_reg (
	.SI(Samples[2]),
	.SE(test_se),
	.RN(RST),
	.Q(sampled_bit),
	.D(N58),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	sampled_bit, 
	Enable, 
	edge_count, 
	Prescale, 
	P_DATA, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input sampled_bit;
   input Enable;
   input [5:0] edge_count;
   input [5:0] Prescale;
   output [7:0] P_DATA;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N1;
   wire N2;
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire n1;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;

   assign test_so = n24 ;

   // Module instantiations
   OAI22X1M U3 (
	.Y(n11),
	.B1(n29),
	.B0(n1),
	.A1(n30),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U4 (
	.Y(n12),
	.B1(n28),
	.B0(n1),
	.A1(n29),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U5 (
	.Y(n13),
	.B1(n27),
	.B0(n1),
	.A1(n28),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U6 (
	.Y(n14),
	.B1(n26),
	.B0(n1),
	.A1(n27),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U7 (
	.Y(n15),
	.B1(n25),
	.B0(n1),
	.A1(n26),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U8 (
	.Y(n16),
	.B1(n24),
	.B0(n1),
	.A1(n25),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n31),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(n1),
	.B(Enable),
	.A(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U11 (
	.Y(n10),
	.B1(n30),
	.B0(n1),
	.A1N(n1),
	.A0N(P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U12 (
	.Y(n17),
	.B1(n24),
	.B0(n31),
	.A1N(n31),
	.A0N(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U13 (
	.Y(n2),
	.B(Prescale[0]),
	.A(Prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n6),
	.A(Prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n29),
	.A(P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n25),
	.A(P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n24),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n28),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n30),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n27),
	.A(P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n26),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U22 (
	.Y(N1),
	.A(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U23 (
	.Y(N2),
	.B0(n2),
	.A1N(Prescale[1]),
	.A0N(Prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(n3),
	.B(Prescale[2]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U25 (
	.Y(N3),
	.B0(n3),
	.A1(Prescale[2]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U26 (
	.Y(n4),
	.B(n6),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U27 (
	.Y(N4),
	.B0(n4),
	.A1(n6),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U28 (
	.Y(N5),
	.B(n4),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U29 (
	.Y(n5),
	.B(n4),
	.A(Prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(N6),
	.B(n5),
	.A(Prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U31 (
	.Y(n7),
	.B(N1),
	.AN(edge_count[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U32 (
	.Y(n19),
	.B1(n7),
	.B0(edge_count[1]),
	.A1N(N2),
	.A0(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U33 (
	.Y(n8),
	.B(edge_count[0]),
	.AN(N1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U34 (
	.Y(n18),
	.B1(n8),
	.B0(N2),
	.A1N(edge_count[1]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U35 (
	.Y(n9),
	.B(edge_count[5]),
	.A(N6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U36 (
	.Y(n23),
	.C(n9),
	.B(n18),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n22),
	.B(edge_count[4]),
	.A(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n21),
	.B(edge_count[2]),
	.A(N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U39 (
	.Y(n20),
	.B(edge_count[3]),
	.A(N4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U40 (
	.Y(N7),
	.D(n20),
	.C(n21),
	.B(n22),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[0]  (
	.SI(sampled_bit),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[0]),
	.D(n10),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[5]  (
	.SI(n27),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[5]),
	.D(n15),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[1]  (
	.SI(P_DATA[0]),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[1]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[4]  (
	.SI(n28),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[4]),
	.D(n14),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[7]  (
	.SI(n25),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[7]),
	.D(n17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[3]  (
	.SI(n29),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[3]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[6]  (
	.SI(n26),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[6]),
	.D(n16),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_reg[2]  (
	.SI(n30),
	.SE(test_se),
	.RN(RST),
	.Q(P_DATA[2]),
	.D(n12),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module strt_chk_test_1 (
	CLK, 
	RST, 
	sampled_bit, 
	Enable, 
	strt_glitch, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input sampled_bit;
   input Enable;
   output strt_glitch;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;

   // Module instantiations
   AO2B2X2M U2 (
	.Y(n1),
	.B1(Enable),
	.B0(sampled_bit),
	.A1N(Enable),
	.A0(strt_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M strt_glitch_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(strt_glitch),
	.D(n1),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module par_chk_DATA_WIDTH8_test_1 (
	CLK, 
	RST, 
	parity_type, 
	sampled_bit, 
	Enable, 
	P_DATA, 
	par_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input parity_type;
   input sampled_bit;
   input Enable;
   input [7:0] P_DATA;
   output par_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n2;
   wire n11;
   wire n12;

   // Module instantiations
   XNOR2X2M U2 (
	.Y(n5),
	.B(parity_type),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U3 (
	.Y(n4),
	.C(n6),
	.B(P_DATA[4]),
	.A(P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(n6),
	.B(P_DATA[6]),
	.A(P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U5 (
	.Y(n3),
	.C(n7),
	.B(P_DATA[0]),
	.A(P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(n7),
	.B(P_DATA[2]),
	.A(P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U7 (
	.Y(n8),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n2),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U9 (
	.Y(n1),
	.C(n5),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U11 (
	.Y(n12),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M par_err_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.QN(n11),
	.Q(par_err),
	.D(n8),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stp_chk_test_1 (
	CLK, 
	RST, 
	sampled_bit, 
	Enable, 
	stp_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input sampled_bit;
   input Enable;
   output stp_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;
   wire n1;
   wire n5;
   wire n6;

   // Module instantiations
   OAI2BB2X1M U2 (
	.Y(n2),
	.B1(n1),
	.B0(sampled_bit),
	.A1N(n1),
	.A0N(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n1),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U5 (
	.Y(n6),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M stp_err_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.QN(n5),
	.Q(stp_err),
	.D(n2),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_CTRL_test_1 (
	clk, 
	rst_n, 
	RX_P_Data, 
	RX_D_VLD, 
	RdData, 
	RdData_Valid, 
	ALU_OUT, 
	OUT_Valid, 
	FIFO_FULL, 
	Address, 
	WrEn, 
	RdEn, 
	WrData, 
	ALU_EN, 
	ALU_FUN, 
	CLK_EN, 
	clk_div_en, 
	WR_DATA, 
	WR_INC, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN2_SYNC_SCAN_RST1, 
	REF_SCAN_CLK__L6_N4, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   input [7:0] RX_P_Data;
   input RX_D_VLD;
   input [7:0] RdData;
   input RdData_Valid;
   input [15:0] ALU_OUT;
   input OUT_Valid;
   input FIFO_FULL;
   output [3:0] Address;
   output WrEn;
   output RdEn;
   output [7:0] WrData;
   output ALU_EN;
   output [3:0] ALU_FUN;
   output CLK_EN;
   output clk_div_en;
   output [7:0] WR_DATA;
   output WR_INC;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN2_SYNC_SCAN_RST1;
   input REF_SCAN_CLK__L6_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire FE_OFN4_Address_3_;
   wire FE_OFN3_Address_2_;
   wire ALU_OUT_BYTE;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n87;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire [3:0] state;

   assign test_so = n13 ;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC4_Address_3_ (
	.Y(Address[3]),
	.A(FE_OFN4_Address_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC3_Address_2_ (
	.Y(Address[2]),
	.A(FE_OFN3_Address_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(ALU_FUN[2]),
	.B(n77),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(ALU_FUN[0]),
	.B(n77),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U7 (
	.Y(FE_OFN3_Address_2_),
	.B1(n25),
	.B0(n71),
	.A1(n16),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2X2M U8 (
	.Y(n27),
	.B1(n8),
	.B0(n3),
	.A1N(RX_D_VLD),
	.A0N(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U9 (
	.Y(n58),
	.B(n55),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n10),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U11 (
	.Y(RdEn),
	.B(n20),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U12 (
	.Y(n55),
	.C(n38),
	.B(n48),
	.A(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U13 (
	.Y(n56),
	.B(n76),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n6),
	.A(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(WrData[0]),
	.B(n58),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(WrData[1]),
	.B(n58),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(WrData[2]),
	.B(n58),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(WrData[3]),
	.B(n58),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(WrData[4]),
	.B(n58),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U20 (
	.Y(WrData[6]),
	.B(n58),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(WrData[7]),
	.B(n58),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U22 (
	.Y(n57),
	.B(n60),
	.AN(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(WR_INC),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U24 (
	.Y(n85),
	.B0(n42),
	.A1(n7),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U25 (
	.Y(n42),
	.B0(n27),
	.A2(n30),
	.A1(n6),
	.A0(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n8),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(WrEn),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U28 (
	.Y(ALU_EN),
	.B(n77),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U29 (
	.Y(n61),
	.B(n3),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n9),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n12),
	.A(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n11),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(ALU_FUN[1]),
	.B(n77),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U34 (
	.Y(ALU_FUN[3]),
	.B(n77),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U35 (
	.Y(CLK_EN),
	.B(n44),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U36 (
	.Y(FE_OFN4_Address_3_),
	.B1(n24),
	.B0(n71),
	.A1(n15),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U37 (
	.Y(Address[0]),
	.C1(n48),
	.C0(n20),
	.B1(n18),
	.B0(n4),
	.A1(n87),
	.A0(n71), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U38 (
	.Y(n71),
	.B0(RdEn),
	.A1(RX_D_VLD),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U39 (
	.Y(n76),
	.B(state[3]),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U40 (
	.Y(Address[1]),
	.B1(n26),
	.B0(n71),
	.A1(n17),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U41 (
	.Y(n51),
	.B(state[3]),
	.A(state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U42 (
	.Y(n52),
	.B(state[1]),
	.A(state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U43 (
	.Y(n75),
	.C(state[1]),
	.B(n7),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U44 (
	.Y(n38),
	.C(state[0]),
	.B(n19),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U45 (
	.Y(n48),
	.C(n76),
	.B(n7),
	.A(state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U46 (
	.Y(n74),
	.C(state[0]),
	.B(n51),
	.A(state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n19),
	.A(state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n7),
	.A(state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n4),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U50 (
	.Y(n72),
	.C0(RX_D_VLD),
	.B0(n74),
	.A1(n73),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U51 (
	.Y(n73),
	.B(n75),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n20),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n14),
	.A(state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U54 (
	.Y(n54),
	.D(n55),
	.C(n10),
	.B(n6),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U55 (
	.Y(n31),
	.C(n13),
	.B(state[2]),
	.AN(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U56 (
	.Y(n63),
	.B(ALU_OUT_BYTE),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U57 (
	.Y(n44),
	.D(n14),
	.C(n19),
	.B(state[0]),
	.A(state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U58 (
	.Y(WrData[5]),
	.B(n58),
	.AN(RX_P_Data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U59 (
	.Y(n30),
	.B0(n45),
	.A1(n44),
	.A0(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U60 (
	.Y(n43),
	.B(FIFO_FULL),
	.AN(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U61 (
	.Y(n83),
	.C0(n32),
	.B0(n5),
	.A1(n14),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U62 (
	.Y(n32),
	.B0(n12),
	.A2(n33),
	.A1(RX_P_Data[4]),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U63 (
	.Y(n5),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U64 (
	.Y(n33),
	.C(RX_P_Data[2]),
	.B(RX_P_Data[6]),
	.A(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U65 (
	.Y(n82),
	.C0(n29),
	.B0(n28),
	.A1(n13),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U66 (
	.Y(n28),
	.B0(n31),
	.A1N(RdData_Valid),
	.A0(FIFO_FULL), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U67 (
	.Y(n29),
	.B0(n27),
	.A1(n30),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U68 (
	.Y(n59),
	.B(n8),
	.A(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U69 (
	.Y(n25),
	.A(RX_P_Data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U70 (
	.Y(n87),
	.A(RX_P_Data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U71 (
	.Y(WR_DATA[0]),
	.B0(n70),
	.A1N(n61),
	.A0N(ALU_OUT[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U72 (
	.Y(n70),
	.B1(n63),
	.B0(ALU_OUT[0]),
	.A1(n60),
	.A0(RdData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U73 (
	.Y(WR_DATA[1]),
	.B0(n69),
	.A1N(n61),
	.A0N(ALU_OUT[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U74 (
	.Y(n69),
	.B1(n63),
	.B0(ALU_OUT[1]),
	.A1(n60),
	.A0(RdData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U75 (
	.Y(WR_DATA[2]),
	.B0(n68),
	.A1N(n61),
	.A0N(ALU_OUT[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U76 (
	.Y(n68),
	.B1(n63),
	.B0(ALU_OUT[2]),
	.A1(n60),
	.A0(RdData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U77 (
	.Y(WR_DATA[3]),
	.B0(n67),
	.A1N(n61),
	.A0N(ALU_OUT[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U78 (
	.Y(n67),
	.B1(n63),
	.B0(ALU_OUT[3]),
	.A1(n60),
	.A0(RdData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U79 (
	.Y(WR_DATA[4]),
	.B0(n66),
	.A1N(n61),
	.A0N(ALU_OUT[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U80 (
	.Y(n66),
	.B1(n63),
	.B0(ALU_OUT[4]),
	.A1(n60),
	.A0(RdData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U81 (
	.Y(WR_DATA[5]),
	.B0(n65),
	.A1N(n61),
	.A0N(ALU_OUT[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U82 (
	.Y(n65),
	.B1(n63),
	.B0(ALU_OUT[5]),
	.A1(n60),
	.A0(RdData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U83 (
	.Y(WR_DATA[6]),
	.B0(n64),
	.A1N(n61),
	.A0N(ALU_OUT[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U84 (
	.Y(n64),
	.B1(n63),
	.B0(ALU_OUT[6]),
	.A1(n60),
	.A0(RdData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U85 (
	.Y(WR_DATA[7]),
	.B0(n62),
	.A1N(n61),
	.A0N(ALU_OUT[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U86 (
	.Y(n62),
	.B1(n63),
	.B0(ALU_OUT[7]),
	.A1(n60),
	.A0(RdData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n80),
	.B1(n17),
	.B0(n6),
	.A1N(n6),
	.A0N(Address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n79),
	.B1(n16),
	.B0(n6),
	.A1N(n6),
	.A0N(Address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n78),
	.B1(n15),
	.B0(n6),
	.A1N(n6),
	.A0N(Address[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n81),
	.B1(n18),
	.B0(n6),
	.A1N(n6),
	.A0N(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U91 (
	.Y(n84),
	.B0(n36),
	.A1(n19),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U92 (
	.Y(n36),
	.B0(n27),
	.A2(n12),
	.A1(n6),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U93 (
	.Y(n37),
	.B0(n40),
	.A2(n34),
	.A1(RX_P_Data[0]),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U94 (
	.Y(n39),
	.C(n25),
	.B(n22),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U95 (
	.Y(n26),
	.A(RX_P_Data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U96 (
	.Y(n60),
	.B(RdData_Valid),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n24),
	.A(RX_P_Data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U98 (
	.Y(n13),
	.A(state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U99 (
	.Y(n86),
	.B1(n3),
	.B0(WR_INC),
	.A2(n57),
	.A1(ALU_OUT_BYTE),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U100 (
	.Y(n41),
	.D(n53),
	.C(n52),
	.B(n51),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U101 (
	.Y(n53),
	.B(n21),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U102 (
	.Y(n45),
	.C(state[0]),
	.B(state[1]),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U103 (
	.Y(n34),
	.C(RX_P_Data[5]),
	.B(RX_P_Data[1]),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U104 (
	.Y(n23),
	.A(RX_P_Data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U105 (
	.Y(n22),
	.A(RX_P_Data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U106 (
	.Y(n35),
	.B(n46),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U107 (
	.Y(n46),
	.D(n47),
	.C(RX_P_Data[6]),
	.B(RX_P_Data[2]),
	.A(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U108 (
	.Y(n47),
	.D(RX_P_Data[0]),
	.C(RX_P_Data[1]),
	.B(RX_P_Data[4]),
	.A(RX_P_Data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U109 (
	.Y(n3),
	.A(ALU_OUT_BYTE), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U110 (
	.Y(n40),
	.B(n49),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U111 (
	.Y(n49),
	.D(n50),
	.C(RX_P_Data[6]),
	.B(n41),
	.A(RX_P_Data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U112 (
	.Y(n50),
	.D(n87),
	.C(n25),
	.B(RX_P_Data[1]),
	.A(RX_P_Data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U113 (
	.Y(n21),
	.A(RX_P_Data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U114 (
	.Y(n77),
	.B(RX_D_VLD),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M ALU_OUT_BYTE_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(ALU_OUT_BYTE),
	.D(n86),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Address_s_reg[0]  (
	.SI(ALU_OUT_BYTE),
	.SE(test_se),
	.RN(rst_n),
	.QN(n18),
	.Q(n93),
	.D(n81),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Address_s_reg[3]  (
	.SI(n91),
	.SE(test_se),
	.RN(rst_n),
	.QN(n15),
	.Q(n92),
	.D(n78),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Address_s_reg[2]  (
	.SI(n90),
	.SE(test_se),
	.RN(rst_n),
	.QN(n16),
	.Q(n91),
	.D(n79),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \Address_s_reg[1]  (
	.SI(n93),
	.SE(test_se),
	.RN(rst_n),
	.QN(n17),
	.Q(n90),
	.D(n80),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \state_reg[2]  (
	.SI(state[1]),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(state[2]),
	.D(n83),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \state_reg[3]  (
	.SI(n14),
	.SE(test_se),
	.RN(FE_OFN2_SYNC_SCAN_RST1),
	.Q(state[3]),
	.D(n82),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \state_reg[0]  (
	.SI(n92),
	.SE(test_se),
	.RN(rst_n),
	.Q(state[0]),
	.D(n85),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \state_reg[1]  (
	.SI(state[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(state[1]),
	.D(n84),
	.CK(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(clk_div_en),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RegFile_WIDTH8_DEPTH16_test_1 (
	CLK, 
	RST, 
	WrEn, 
	RdEn, 
	Address, 
	WrData, 
	RdData, 
	RdData_VLD, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN0_SYNC_SCAN_RST1, 
	FE_OFN1_SYNC_SCAN_RST1, 
	REF_SCAN_CLK__L6_N1, 
	REF_SCAN_CLK__L6_N10, 
	REF_SCAN_CLK__L6_N11, 
	REF_SCAN_CLK__L6_N2, 
	REF_SCAN_CLK__L6_N3, 
	REF_SCAN_CLK__L6_N7, 
	REF_SCAN_CLK__L6_N8, 
	REF_SCAN_CLK__L6_N9, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input WrEn;
   input RdEn;
   input [3:0] Address;
   input [7:0] WrData;
   output [7:0] RdData;
   output RdData_VLD;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN0_SYNC_SCAN_RST1;
   input FE_OFN1_SYNC_SCAN_RST1;
   input REF_SCAN_CLK__L6_N1;
   input REF_SCAN_CLK__L6_N10;
   input REF_SCAN_CLK__L6_N11;
   input REF_SCAN_CLK__L6_N2;
   input REF_SCAN_CLK__L6_N3;
   input REF_SCAN_CLK__L6_N7;
   input REF_SCAN_CLK__L6_N8;
   input REF_SCAN_CLK__L6_N9;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN6_SO_1_;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire \regArr[15][7] ;
   wire \regArr[15][6] ;
   wire \regArr[15][5] ;
   wire \regArr[15][4] ;
   wire \regArr[15][3] ;
   wire \regArr[15][2] ;
   wire \regArr[15][1] ;
   wire \regArr[15][0] ;
   wire \regArr[14][7] ;
   wire \regArr[14][6] ;
   wire \regArr[14][5] ;
   wire \regArr[14][4] ;
   wire \regArr[14][3] ;
   wire \regArr[14][2] ;
   wire \regArr[14][1] ;
   wire \regArr[14][0] ;
   wire \regArr[13][7] ;
   wire \regArr[13][6] ;
   wire \regArr[13][5] ;
   wire \regArr[13][4] ;
   wire \regArr[13][3] ;
   wire \regArr[13][2] ;
   wire \regArr[13][1] ;
   wire \regArr[13][0] ;
   wire \regArr[12][7] ;
   wire \regArr[12][6] ;
   wire \regArr[12][5] ;
   wire \regArr[12][4] ;
   wire \regArr[12][3] ;
   wire \regArr[12][2] ;
   wire \regArr[12][1] ;
   wire \regArr[12][0] ;
   wire \regArr[11][7] ;
   wire \regArr[11][6] ;
   wire \regArr[11][5] ;
   wire \regArr[11][4] ;
   wire \regArr[11][3] ;
   wire \regArr[11][2] ;
   wire \regArr[11][1] ;
   wire \regArr[11][0] ;
   wire \regArr[10][7] ;
   wire \regArr[10][6] ;
   wire \regArr[10][5] ;
   wire \regArr[10][4] ;
   wire \regArr[10][3] ;
   wire \regArr[10][2] ;
   wire \regArr[10][1] ;
   wire \regArr[10][0] ;
   wire \regArr[9][7] ;
   wire \regArr[9][6] ;
   wire \regArr[9][5] ;
   wire \regArr[9][4] ;
   wire \regArr[9][3] ;
   wire \regArr[9][2] ;
   wire \regArr[9][1] ;
   wire \regArr[9][0] ;
   wire \regArr[8][7] ;
   wire \regArr[8][6] ;
   wire \regArr[8][5] ;
   wire \regArr[8][4] ;
   wire \regArr[8][3] ;
   wire \regArr[8][2] ;
   wire \regArr[8][1] ;
   wire \regArr[8][0] ;
   wire \regArr[7][7] ;
   wire \regArr[7][6] ;
   wire \regArr[7][5] ;
   wire \regArr[7][4] ;
   wire \regArr[7][3] ;
   wire \regArr[7][2] ;
   wire \regArr[7][1] ;
   wire \regArr[7][0] ;
   wire \regArr[6][7] ;
   wire \regArr[6][6] ;
   wire \regArr[6][5] ;
   wire \regArr[6][4] ;
   wire \regArr[6][3] ;
   wire \regArr[6][2] ;
   wire \regArr[6][1] ;
   wire \regArr[6][0] ;
   wire \regArr[5][7] ;
   wire \regArr[5][6] ;
   wire \regArr[5][5] ;
   wire \regArr[5][4] ;
   wire \regArr[5][3] ;
   wire \regArr[5][2] ;
   wire \regArr[5][1] ;
   wire \regArr[5][0] ;
   wire \regArr[4][7] ;
   wire \regArr[4][6] ;
   wire \regArr[4][5] ;
   wire \regArr[4][4] ;
   wire \regArr[4][3] ;
   wire \regArr[4][2] ;
   wire \regArr[4][1] ;
   wire \regArr[4][0] ;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n199;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n242;
   wire n229;

   assign N11 = Address[0] ;
   assign N12 = Address[1] ;
   assign N13 = Address[2] ;
   assign N14 = Address[3] ;
   assign test_so2 = \regArr[15][7]  ;
   assign test_so1 = \regArr[13][4]  ;

   // Module instantiations
   BUFX10M FE_OFC6_SO_1_ (
	.Y(\regArr[13][4] ),
	.A(FE_OFN6_SO_1_), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U3 (
	.Y(n23),
	.B(n199),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(n26),
	.B(n204),
	.AN(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U5 (
	.Y(n20),
	.B(N13),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n15),
	.B(N13),
	.A(n199), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U7 (
	.Y(n201),
	.A(n203), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n199),
	.A(n204), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U10 (
	.Y(n202),
	.A(n203), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n228),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U13 (
	.Y(n30),
	.B(N11),
	.AN(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U14 (
	.Y(n32),
	.B(n203),
	.AN(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U15 (
	.Y(n29),
	.B(n15),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(n31),
	.B(n15),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U17 (
	.Y(n33),
	.B(n20),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n34),
	.B(n20),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(n35),
	.B(n23),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U20 (
	.Y(n36),
	.B(n23),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U21 (
	.Y(n37),
	.B(n26),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(n39),
	.B(n26),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U23 (
	.Y(n16),
	.B(N11),
	.AN(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U24 (
	.Y(n18),
	.B(n203),
	.AN(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(n17),
	.B(n15),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U26 (
	.Y(n19),
	.B(n16),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U27 (
	.Y(n21),
	.B(n18),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U28 (
	.Y(n22),
	.B(n16),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U29 (
	.Y(n24),
	.B(n18),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U30 (
	.Y(n25),
	.B(n16),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U31 (
	.Y(n28),
	.B(n18),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n14),
	.B(n16),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U33 (
	.Y(n12),
	.B(RdEn),
	.AN(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U34 (
	.Y(n13),
	.B(RdEn),
	.AN(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U45 (
	.Y(n38),
	.B(n13),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n203),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n204),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n220),
	.A(WrData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n221),
	.A(WrData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n222),
	.A(WrData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U51 (
	.Y(n223),
	.A(WrData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n224),
	.A(WrData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n226),
	.A(WrData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U54 (
	.Y(n227),
	.A(WrData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U55 (
	.Y(n27),
	.B(N14),
	.AN(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U61 (
	.Y(n113),
	.B1(n29),
	.B0(n220),
	.A1N(n29),
	.A0N(\regArr[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U62 (
	.Y(n114),
	.B1(n29),
	.B0(n221),
	.A1N(n29),
	.A0N(\regArr[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U63 (
	.Y(n115),
	.B1(n29),
	.B0(n222),
	.A1N(n29),
	.A0N(\regArr[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U64 (
	.Y(n116),
	.B1(n29),
	.B0(n223),
	.A1N(n29),
	.A0N(\regArr[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U65 (
	.Y(n117),
	.B1(n29),
	.B0(n224),
	.A1N(n29),
	.A0N(\regArr[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U66 (
	.Y(n118),
	.B1(n29),
	.B0(n225),
	.A1N(n29),
	.A0N(\regArr[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U67 (
	.Y(n119),
	.B1(n29),
	.B0(n226),
	.A1N(n29),
	.A0N(\regArr[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U68 (
	.Y(n120),
	.B1(n29),
	.B0(n227),
	.A1N(n29),
	.A0N(\regArr[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U69 (
	.Y(n121),
	.B1(n31),
	.B0(n220),
	.A1N(n31),
	.A0N(\regArr[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U70 (
	.Y(n122),
	.B1(n31),
	.B0(n221),
	.A1N(n31),
	.A0N(\regArr[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U71 (
	.Y(n123),
	.B1(n31),
	.B0(n222),
	.A1N(n31),
	.A0N(\regArr[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U72 (
	.Y(n124),
	.B1(n31),
	.B0(n223),
	.A1N(n31),
	.A0N(\regArr[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U73 (
	.Y(n125),
	.B1(n31),
	.B0(n224),
	.A1N(n31),
	.A0N(\regArr[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U74 (
	.Y(n126),
	.B1(n31),
	.B0(n225),
	.A1N(n31),
	.A0N(\regArr[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U75 (
	.Y(n127),
	.B1(n31),
	.B0(n226),
	.A1N(n31),
	.A0N(\regArr[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U76 (
	.Y(n128),
	.B1(n31),
	.B0(n227),
	.A1N(n31),
	.A0N(\regArr[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U77 (
	.Y(n129),
	.B1(n33),
	.B0(n220),
	.A1N(n33),
	.A0N(\regArr[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U78 (
	.Y(n130),
	.B1(n33),
	.B0(n221),
	.A1N(n33),
	.A0N(\regArr[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U79 (
	.Y(n131),
	.B1(n33),
	.B0(n222),
	.A1N(n33),
	.A0N(\regArr[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U80 (
	.Y(n132),
	.B1(n33),
	.B0(n223),
	.A1N(n33),
	.A0N(\regArr[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U81 (
	.Y(n133),
	.B1(n33),
	.B0(n224),
	.A1N(n33),
	.A0N(\regArr[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U82 (
	.Y(n134),
	.B1(n33),
	.B0(n225),
	.A1N(n33),
	.A0N(\regArr[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U83 (
	.Y(n135),
	.B1(n33),
	.B0(n226),
	.A1N(n33),
	.A0N(\regArr[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n136),
	.B1(n33),
	.B0(n227),
	.A1N(n33),
	.A0N(\regArr[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n137),
	.B1(n34),
	.B0(n220),
	.A1N(n34),
	.A0N(\regArr[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n138),
	.B1(n34),
	.B0(n221),
	.A1N(n34),
	.A0N(\regArr[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n139),
	.B1(n34),
	.B0(n222),
	.A1N(n34),
	.A0N(\regArr[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n140),
	.B1(n34),
	.B0(n223),
	.A1N(n34),
	.A0N(\regArr[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n141),
	.B1(n34),
	.B0(n224),
	.A1N(n34),
	.A0N(\regArr[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n142),
	.B1(n34),
	.B0(n225),
	.A1N(n34),
	.A0N(\regArr[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n143),
	.B1(n34),
	.B0(n226),
	.A1N(n34),
	.A0N(\regArr[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U92 (
	.Y(n144),
	.B1(n34),
	.B0(n227),
	.A1N(n34),
	.A0N(\regArr[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U93 (
	.Y(n145),
	.B1(n35),
	.B0(n220),
	.A1N(n35),
	.A0N(\regArr[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U94 (
	.Y(n146),
	.B1(n35),
	.B0(n221),
	.A1N(n35),
	.A0N(\regArr[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n147),
	.B1(n35),
	.B0(n222),
	.A1N(n35),
	.A0N(\regArr[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U96 (
	.Y(n148),
	.B1(n35),
	.B0(n223),
	.A1N(n35),
	.A0N(\regArr[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U97 (
	.Y(n149),
	.B1(n35),
	.B0(n224),
	.A1N(n35),
	.A0N(\regArr[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U98 (
	.Y(n150),
	.B1(n35),
	.B0(n225),
	.A1N(n35),
	.A0N(\regArr[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U99 (
	.Y(n151),
	.B1(n35),
	.B0(n226),
	.A1N(n35),
	.A0N(\regArr[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n152),
	.B1(n35),
	.B0(n227),
	.A1N(n35),
	.A0N(\regArr[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n153),
	.B1(n36),
	.B0(n220),
	.A1N(n36),
	.A0N(\regArr[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n154),
	.B1(n36),
	.B0(n221),
	.A1N(n36),
	.A0N(\regArr[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n155),
	.B1(n36),
	.B0(n222),
	.A1N(n36),
	.A0N(\regArr[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n156),
	.B1(n36),
	.B0(n223),
	.A1N(n36),
	.A0N(\regArr[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U105 (
	.Y(n157),
	.B1(n36),
	.B0(n224),
	.A1N(n36),
	.A0N(n240), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U106 (
	.Y(n158),
	.B1(n36),
	.B0(n225),
	.A1N(n36),
	.A0N(\regArr[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U107 (
	.Y(n159),
	.B1(n36),
	.B0(n226),
	.A1N(n36),
	.A0N(\regArr[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U108 (
	.Y(n160),
	.B1(n36),
	.B0(n227),
	.A1N(n36),
	.A0N(\regArr[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U109 (
	.Y(n161),
	.B1(n37),
	.B0(n220),
	.A1N(n37),
	.A0N(\regArr[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U110 (
	.Y(n162),
	.B1(n37),
	.B0(n221),
	.A1N(n37),
	.A0N(\regArr[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U111 (
	.Y(n163),
	.B1(n37),
	.B0(n222),
	.A1N(n37),
	.A0N(\regArr[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U112 (
	.Y(n164),
	.B1(n37),
	.B0(n223),
	.A1N(n37),
	.A0N(\regArr[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U113 (
	.Y(n165),
	.B1(n37),
	.B0(n224),
	.A1N(n37),
	.A0N(\regArr[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U114 (
	.Y(n166),
	.B1(n37),
	.B0(n225),
	.A1N(n37),
	.A0N(\regArr[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U115 (
	.Y(n167),
	.B1(n37),
	.B0(n226),
	.A1N(n37),
	.A0N(\regArr[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U116 (
	.Y(n168),
	.B1(n37),
	.B0(n227),
	.A1N(n37),
	.A0N(\regArr[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U117 (
	.Y(n169),
	.B1(n39),
	.B0(n220),
	.A1N(n39),
	.A0N(\regArr[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n170),
	.B1(n39),
	.B0(n221),
	.A1N(n39),
	.A0N(\regArr[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n171),
	.B1(n39),
	.B0(n222),
	.A1N(n39),
	.A0N(\regArr[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n172),
	.B1(n39),
	.B0(n223),
	.A1N(n39),
	.A0N(\regArr[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n173),
	.B1(n39),
	.B0(n224),
	.A1N(n39),
	.A0N(\regArr[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n174),
	.B1(n39),
	.B0(n225),
	.A1N(n39),
	.A0N(\regArr[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n175),
	.B1(n39),
	.B0(n226),
	.A1N(n39),
	.A0N(\regArr[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n176),
	.B1(n39),
	.B0(n227),
	.A1N(n39),
	.A0N(\regArr[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U125 (
	.Y(n40),
	.B1(n12),
	.B0(RdData[0]),
	.A1(n228),
	.A0(N43), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U126 (
	.Y(N43),
	.S1(N13),
	.S0(N14),
	.D(n1),
	.C(n3),
	.B(n2),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U127 (
	.Y(n4),
	.S1(n199),
	.S0(N11),
	.D(REG3[0]),
	.C(REG2[0]),
	.B(REG1[0]),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U128 (
	.Y(n2),
	.S1(n199),
	.S0(N11),
	.D(\regArr[11][0] ),
	.C(\regArr[10][0] ),
	.B(\regArr[9][0] ),
	.A(\regArr[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U129 (
	.Y(n41),
	.B1(n12),
	.B0(RdData[1]),
	.A1(n228),
	.A0(N42), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U130 (
	.Y(N42),
	.S1(N13),
	.S0(N14),
	.D(n5),
	.C(n7),
	.B(n6),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U131 (
	.Y(n6),
	.S1(n199),
	.S0(N11),
	.D(\regArr[11][1] ),
	.C(\regArr[10][1] ),
	.B(\regArr[9][1] ),
	.A(\regArr[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U132 (
	.Y(n5),
	.S1(n199),
	.S0(n201),
	.D(\regArr[15][1] ),
	.C(\regArr[14][1] ),
	.B(\regArr[13][1] ),
	.A(\regArr[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U133 (
	.Y(n42),
	.B1(n12),
	.B0(RdData[2]),
	.A1(n228),
	.A0(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U134 (
	.Y(N41),
	.S1(N13),
	.S0(N14),
	.D(n9),
	.C(n11),
	.B(n10),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U135 (
	.Y(n177),
	.S1(N12),
	.S0(n201),
	.D(REG3[2]),
	.C(REG2[2]),
	.B(REG1[2]),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U136 (
	.Y(n10),
	.S1(N12),
	.S0(n201),
	.D(\regArr[11][2] ),
	.C(\regArr[10][2] ),
	.B(\regArr[9][2] ),
	.A(\regArr[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U137 (
	.Y(n43),
	.B1(n12),
	.B0(RdData[3]),
	.A1(n228),
	.A0(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U138 (
	.Y(N40),
	.S1(N13),
	.S0(N14),
	.D(n178),
	.C(n180),
	.B(n179),
	.A(n181), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U139 (
	.Y(n181),
	.S1(N12),
	.S0(n201),
	.D(REG3[3]),
	.C(REG2[3]),
	.B(REG1[3]),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U140 (
	.Y(n179),
	.S1(N12),
	.S0(n201),
	.D(\regArr[11][3] ),
	.C(\regArr[10][3] ),
	.B(\regArr[9][3] ),
	.A(\regArr[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U141 (
	.Y(n44),
	.B1(n12),
	.B0(RdData[4]),
	.A1(n228),
	.A0(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U142 (
	.Y(N39),
	.S1(N13),
	.S0(N14),
	.D(n182),
	.C(n184),
	.B(n183),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U143 (
	.Y(n185),
	.S1(N12),
	.S0(n202),
	.D(REG3[4]),
	.C(REG2[4]),
	.B(REG1[4]),
	.A(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U144 (
	.Y(n183),
	.S1(N12),
	.S0(n201),
	.D(\regArr[11][4] ),
	.C(\regArr[10][4] ),
	.B(\regArr[9][4] ),
	.A(\regArr[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U145 (
	.Y(n45),
	.B1(n12),
	.B0(RdData[5]),
	.A1(n228),
	.A0(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U146 (
	.Y(N38),
	.S1(N13),
	.S0(N14),
	.D(n186),
	.C(n188),
	.B(n187),
	.A(n189), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U147 (
	.Y(n189),
	.S1(N12),
	.S0(n202),
	.D(REG3[5]),
	.C(REG2[5]),
	.B(REG1[5]),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U148 (
	.Y(n187),
	.S1(N12),
	.S0(n202),
	.D(\regArr[11][5] ),
	.C(\regArr[10][5] ),
	.B(\regArr[9][5] ),
	.A(\regArr[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U149 (
	.Y(n46),
	.B1(n12),
	.B0(RdData[6]),
	.A1(n228),
	.A0(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U150 (
	.Y(N37),
	.S1(N13),
	.S0(N14),
	.D(n190),
	.C(n192),
	.B(n191),
	.A(n193), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U151 (
	.Y(n193),
	.S1(N12),
	.S0(n202),
	.D(REG3[6]),
	.C(REG2[6]),
	.B(REG1[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U152 (
	.Y(n191),
	.S1(N12),
	.S0(n202),
	.D(\regArr[11][6] ),
	.C(\regArr[10][6] ),
	.B(\regArr[9][6] ),
	.A(\regArr[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U153 (
	.Y(n47),
	.B1(n12),
	.B0(RdData[7]),
	.A1(n228),
	.A0(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U154 (
	.Y(N36),
	.S1(N13),
	.S0(N14),
	.D(n194),
	.C(n196),
	.B(n195),
	.A(n197), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U155 (
	.Y(n197),
	.S1(N12),
	.S0(n202),
	.D(REG3[7]),
	.C(REG2[7]),
	.B(REG1[7]),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U156 (
	.Y(n195),
	.S1(N12),
	.S0(n202),
	.D(\regArr[11][7] ),
	.C(\regArr[10][7] ),
	.B(\regArr[9][7] ),
	.A(\regArr[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U157 (
	.Y(n8),
	.S1(n199),
	.S0(n201),
	.D(REG3[1]),
	.C(REG2[1]),
	.B(REG1[1]),
	.A(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U158 (
	.Y(n3),
	.S1(n199),
	.S0(N11),
	.D(\regArr[7][0] ),
	.C(\regArr[6][0] ),
	.B(\regArr[5][0] ),
	.A(\regArr[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U159 (
	.Y(n7),
	.S1(n199),
	.S0(n201),
	.D(\regArr[7][1] ),
	.C(\regArr[6][1] ),
	.B(\regArr[5][1] ),
	.A(\regArr[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U160 (
	.Y(n11),
	.S1(N12),
	.S0(n201),
	.D(\regArr[7][2] ),
	.C(\regArr[6][2] ),
	.B(\regArr[5][2] ),
	.A(\regArr[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U161 (
	.Y(n180),
	.S1(N12),
	.S0(n201),
	.D(\regArr[7][3] ),
	.C(\regArr[6][3] ),
	.B(\regArr[5][3] ),
	.A(\regArr[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U162 (
	.Y(n184),
	.S1(N12),
	.S0(n201),
	.D(\regArr[7][4] ),
	.C(\regArr[6][4] ),
	.B(\regArr[5][4] ),
	.A(\regArr[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U163 (
	.Y(n188),
	.S1(N12),
	.S0(n202),
	.D(\regArr[7][5] ),
	.C(\regArr[6][5] ),
	.B(\regArr[5][5] ),
	.A(\regArr[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U164 (
	.Y(n192),
	.S1(N12),
	.S0(n202),
	.D(\regArr[7][6] ),
	.C(\regArr[6][6] ),
	.B(\regArr[5][6] ),
	.A(\regArr[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U165 (
	.Y(n196),
	.S1(N12),
	.S0(n202),
	.D(\regArr[7][7] ),
	.C(\regArr[6][7] ),
	.B(\regArr[5][7] ),
	.A(\regArr[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U166 (
	.Y(n1),
	.S1(n199),
	.S0(n202),
	.D(\regArr[15][0] ),
	.C(\regArr[14][0] ),
	.B(\regArr[13][0] ),
	.A(\regArr[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U167 (
	.Y(n9),
	.S1(n199),
	.S0(n201),
	.D(\regArr[15][2] ),
	.C(\regArr[14][2] ),
	.B(\regArr[13][2] ),
	.A(\regArr[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U168 (
	.Y(n178),
	.S1(n199),
	.S0(n201),
	.D(\regArr[15][3] ),
	.C(\regArr[14][3] ),
	.B(\regArr[13][3] ),
	.A(\regArr[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U169 (
	.Y(n182),
	.S1(N12),
	.S0(n201),
	.D(\regArr[15][4] ),
	.C(\regArr[14][4] ),
	.B(n240),
	.A(\regArr[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U170 (
	.Y(n186),
	.S1(n199),
	.S0(n202),
	.D(\regArr[15][5] ),
	.C(\regArr[14][5] ),
	.B(\regArr[13][5] ),
	.A(\regArr[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U171 (
	.Y(n190),
	.S1(n199),
	.S0(n202),
	.D(\regArr[15][6] ),
	.C(\regArr[14][6] ),
	.B(\regArr[13][6] ),
	.A(\regArr[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U172 (
	.Y(n194),
	.S1(n199),
	.S0(n202),
	.D(\regArr[15][7] ),
	.C(\regArr[14][7] ),
	.B(\regArr[13][7] ),
	.A(\regArr[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U173 (
	.Y(n225),
	.A(WrData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U174 (
	.Y(n49),
	.B1(n220),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U175 (
	.Y(n50),
	.B1(n221),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U176 (
	.Y(n51),
	.B1(n222),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U177 (
	.Y(n52),
	.B1(n223),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U178 (
	.Y(n53),
	.B1(n224),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U179 (
	.Y(n54),
	.B1(n225),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U180 (
	.Y(n55),
	.B1(n226),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U181 (
	.Y(n56),
	.B1(n227),
	.B0(n14),
	.A1N(n14),
	.A0N(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U182 (
	.Y(n57),
	.B1(n17),
	.B0(n220),
	.A1N(n17),
	.A0N(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U183 (
	.Y(n58),
	.B1(n17),
	.B0(n221),
	.A1N(n17),
	.A0N(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U184 (
	.Y(n59),
	.B1(n17),
	.B0(n222),
	.A1N(n17),
	.A0N(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U185 (
	.Y(n60),
	.B1(n17),
	.B0(n223),
	.A1N(n17),
	.A0N(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U186 (
	.Y(n61),
	.B1(n17),
	.B0(n224),
	.A1N(n17),
	.A0N(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U187 (
	.Y(n62),
	.B1(n17),
	.B0(n225),
	.A1N(n17),
	.A0N(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U188 (
	.Y(n63),
	.B1(n17),
	.B0(n226),
	.A1N(n17),
	.A0N(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U189 (
	.Y(n64),
	.B1(n17),
	.B0(n227),
	.A1N(n17),
	.A0N(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U190 (
	.Y(n81),
	.B1(n22),
	.B0(n220),
	.A1N(n22),
	.A0N(\regArr[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U191 (
	.Y(n82),
	.B1(n22),
	.B0(n221),
	.A1N(n22),
	.A0N(\regArr[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U192 (
	.Y(n83),
	.B1(n22),
	.B0(n222),
	.A1N(n22),
	.A0N(\regArr[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U193 (
	.Y(n84),
	.B1(n22),
	.B0(n223),
	.A1N(n22),
	.A0N(\regArr[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U194 (
	.Y(n85),
	.B1(n22),
	.B0(n224),
	.A1N(n22),
	.A0N(\regArr[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U195 (
	.Y(n86),
	.B1(n22),
	.B0(n225),
	.A1N(n22),
	.A0N(\regArr[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U196 (
	.Y(n87),
	.B1(n22),
	.B0(n226),
	.A1N(n22),
	.A0N(\regArr[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U197 (
	.Y(n88),
	.B1(n22),
	.B0(n227),
	.A1N(n22),
	.A0N(\regArr[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U198 (
	.Y(n89),
	.B1(n24),
	.B0(n220),
	.A1N(n24),
	.A0N(\regArr[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U199 (
	.Y(n90),
	.B1(n24),
	.B0(n221),
	.A1N(n24),
	.A0N(\regArr[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U200 (
	.Y(n91),
	.B1(n24),
	.B0(n222),
	.A1N(n24),
	.A0N(\regArr[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U201 (
	.Y(n92),
	.B1(n24),
	.B0(n223),
	.A1N(n24),
	.A0N(\regArr[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U202 (
	.Y(n93),
	.B1(n24),
	.B0(n224),
	.A1N(n24),
	.A0N(\regArr[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U203 (
	.Y(n94),
	.B1(n24),
	.B0(n225),
	.A1N(n24),
	.A0N(\regArr[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U204 (
	.Y(n95),
	.B1(n24),
	.B0(n226),
	.A1N(n24),
	.A0N(\regArr[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U205 (
	.Y(n96),
	.B1(n24),
	.B0(n227),
	.A1N(n24),
	.A0N(\regArr[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U206 (
	.Y(n97),
	.B1(n25),
	.B0(n220),
	.A1N(n25),
	.A0N(\regArr[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n98),
	.B1(n25),
	.B0(n221),
	.A1N(n25),
	.A0N(\regArr[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n99),
	.B1(n25),
	.B0(n222),
	.A1N(n25),
	.A0N(\regArr[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n100),
	.B1(n25),
	.B0(n223),
	.A1N(n25),
	.A0N(\regArr[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n101),
	.B1(n25),
	.B0(n224),
	.A1N(n25),
	.A0N(\regArr[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n102),
	.B1(n25),
	.B0(n225),
	.A1N(n25),
	.A0N(\regArr[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n103),
	.B1(n25),
	.B0(n226),
	.A1N(n25),
	.A0N(\regArr[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n104),
	.B1(n25),
	.B0(n227),
	.A1N(n25),
	.A0N(\regArr[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n105),
	.B1(n28),
	.B0(n220),
	.A1N(n28),
	.A0N(\regArr[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n106),
	.B1(n28),
	.B0(n221),
	.A1N(n28),
	.A0N(\regArr[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n107),
	.B1(n28),
	.B0(n222),
	.A1N(n28),
	.A0N(\regArr[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n108),
	.B1(n28),
	.B0(n223),
	.A1N(n28),
	.A0N(\regArr[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n109),
	.B1(n28),
	.B0(n224),
	.A1N(n28),
	.A0N(\regArr[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n110),
	.B1(n28),
	.B0(n225),
	.A1N(n28),
	.A0N(\regArr[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n111),
	.B1(n28),
	.B0(n226),
	.A1N(n28),
	.A0N(\regArr[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n112),
	.B1(n28),
	.B0(n227),
	.A1N(n28),
	.A0N(\regArr[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n66),
	.B1(n19),
	.B0(n221),
	.A1N(n19),
	.A0N(REG2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n67),
	.B1(n19),
	.B0(n222),
	.A1N(n19),
	.A0N(REG2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n68),
	.B1(n19),
	.B0(n223),
	.A1N(n19),
	.A0N(REG2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n69),
	.B1(n19),
	.B0(n224),
	.A1N(n19),
	.A0N(REG2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n70),
	.B1(n19),
	.B0(n225),
	.A1N(n19),
	.A0N(REG2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n71),
	.B1(n19),
	.B0(n226),
	.A1N(n19),
	.A0N(REG2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n73),
	.B1(n21),
	.B0(n220),
	.A1N(n21),
	.A0N(REG3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n74),
	.B1(n21),
	.B0(n221),
	.A1N(n21),
	.A0N(REG3[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n75),
	.B1(n21),
	.B0(n222),
	.A1N(n21),
	.A0N(REG3[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n76),
	.B1(n21),
	.B0(n223),
	.A1N(n21),
	.A0N(REG3[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n77),
	.B1(n21),
	.B0(n224),
	.A1N(n21),
	.A0N(REG3[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n79),
	.B1(n21),
	.B0(n226),
	.A1N(n21),
	.A0N(REG3[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n80),
	.B1(n21),
	.B0(n227),
	.A1N(n21),
	.A0N(REG3[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n65),
	.B1(n19),
	.B0(n220),
	.A1N(n19),
	.A0N(REG2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n72),
	.B1(n19),
	.B0(n227),
	.A1N(n19),
	.A0N(REG2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n78),
	.B1(n21),
	.B0(n225),
	.A1N(n21),
	.A0N(REG3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U238 (
	.Y(n48),
	.B0(n12),
	.A1N(n13),
	.A0N(RdData_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][7]  (
	.SI(\regArr[13][6] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[13][7] ),
	.D(n160),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][6]  (
	.SI(\regArr[13][5] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[13][6] ),
	.D(n159),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][5]  (
	.SI(test_si3),
	.SE(n234),
	.RN(RST),
	.Q(\regArr[13][5] ),
	.D(n158),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][3]  (
	.SI(\regArr[13][2] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[13][3] ),
	.D(n156),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][2]  (
	.SI(\regArr[13][1] ),
	.SE(n233),
	.RN(RST),
	.Q(\regArr[13][2] ),
	.D(n155),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][1]  (
	.SI(\regArr[13][0] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[13][1] ),
	.D(n154),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[13][0]  (
	.SI(\regArr[12][7] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[13][0] ),
	.D(n153),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][7]  (
	.SI(\regArr[9][6] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][7] ),
	.D(n128),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][6]  (
	.SI(\regArr[9][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][6] ),
	.D(n127),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][5]  (
	.SI(\regArr[9][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][5] ),
	.D(n126),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][4]  (
	.SI(\regArr[9][3] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][4] ),
	.D(n125),
	.CK(REF_SCAN_CLK__L6_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][3]  (
	.SI(\regArr[9][2] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][3] ),
	.D(n124),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][2]  (
	.SI(\regArr[9][1] ),
	.SE(n233),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][2] ),
	.D(n123),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][1]  (
	.SI(\regArr[9][0] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][1] ),
	.D(n122),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[9][0]  (
	.SI(\regArr[8][7] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[9][0] ),
	.D(n121),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][7]  (
	.SI(\regArr[5][6] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[5][7] ),
	.D(n96),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][6]  (
	.SI(\regArr[5][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[5][6] ),
	.D(n95),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][5]  (
	.SI(\regArr[5][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[5][5] ),
	.D(n94),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][4]  (
	.SI(\regArr[5][3] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[5][4] ),
	.D(n93),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][3]  (
	.SI(\regArr[5][2] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[5][3] ),
	.D(n92),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][2]  (
	.SI(\regArr[5][1] ),
	.SE(n233),
	.RN(RST),
	.Q(\regArr[5][2] ),
	.D(n91),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][1]  (
	.SI(\regArr[5][0] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[5][1] ),
	.D(n90),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[5][0]  (
	.SI(\regArr[4][7] ),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[5][0] ),
	.D(n89),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][7]  (
	.SI(\regArr[15][6] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[15][7] ),
	.D(n176),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][6]  (
	.SI(\regArr[15][5] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[15][6] ),
	.D(n175),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][5]  (
	.SI(\regArr[15][4] ),
	.SE(n234),
	.RN(RST),
	.Q(\regArr[15][5] ),
	.D(n174),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][4]  (
	.SI(\regArr[15][3] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[15][4] ),
	.D(n173),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][3]  (
	.SI(\regArr[15][2] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[15][3] ),
	.D(n172),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][2]  (
	.SI(\regArr[15][1] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[15][2] ),
	.D(n171),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][1]  (
	.SI(\regArr[15][0] ),
	.SE(n233),
	.RN(RST),
	.Q(\regArr[15][1] ),
	.D(n170),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[15][0]  (
	.SI(\regArr[14][7] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[15][0] ),
	.D(n169),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][7]  (
	.SI(\regArr[11][6] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][7] ),
	.D(n144),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][6]  (
	.SI(\regArr[11][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][6] ),
	.D(n143),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][5]  (
	.SI(\regArr[11][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][5] ),
	.D(n142),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][4]  (
	.SI(\regArr[11][3] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][4] ),
	.D(n141),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][3]  (
	.SI(\regArr[11][2] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][3] ),
	.D(n140),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][2]  (
	.SI(\regArr[11][1] ),
	.SE(n233),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][2] ),
	.D(n139),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][1]  (
	.SI(\regArr[11][0] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[11][1] ),
	.D(n138),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[11][0]  (
	.SI(\regArr[10][7] ),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[11][0] ),
	.D(n137),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][7]  (
	.SI(\regArr[7][6] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[7][7] ),
	.D(n112),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][6]  (
	.SI(\regArr[7][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[7][6] ),
	.D(n111),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][5]  (
	.SI(\regArr[7][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[7][5] ),
	.D(n110),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][4]  (
	.SI(\regArr[7][3] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[7][4] ),
	.D(n109),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][3]  (
	.SI(\regArr[7][2] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[7][3] ),
	.D(n108),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][2]  (
	.SI(\regArr[7][1] ),
	.SE(n233),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[7][2] ),
	.D(n107),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][1]  (
	.SI(\regArr[7][0] ),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[7][1] ),
	.D(n106),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[7][0]  (
	.SI(\regArr[6][7] ),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[7][0] ),
	.D(n105),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][7]  (
	.SI(\regArr[14][6] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[14][7] ),
	.D(n168),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][6]  (
	.SI(\regArr[14][5] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[14][6] ),
	.D(n167),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][5]  (
	.SI(\regArr[14][4] ),
	.SE(n234),
	.RN(RST),
	.Q(\regArr[14][5] ),
	.D(n166),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][4]  (
	.SI(\regArr[14][3] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[14][4] ),
	.D(n165),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][3]  (
	.SI(\regArr[14][2] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[14][3] ),
	.D(n164),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][2]  (
	.SI(\regArr[14][1] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[14][2] ),
	.D(n163),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][1]  (
	.SI(\regArr[14][0] ),
	.SE(n233),
	.RN(RST),
	.Q(\regArr[14][1] ),
	.D(n162),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[14][0]  (
	.SI(\regArr[13][7] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[14][0] ),
	.D(n161),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][7]  (
	.SI(\regArr[10][6] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][7] ),
	.D(n136),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][6]  (
	.SI(\regArr[10][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][6] ),
	.D(n135),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][5]  (
	.SI(\regArr[10][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][5] ),
	.D(n134),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][4]  (
	.SI(\regArr[10][3] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][4] ),
	.D(n133),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][3]  (
	.SI(\regArr[10][2] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][3] ),
	.D(n132),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][2]  (
	.SI(\regArr[10][1] ),
	.SE(n233),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][2] ),
	.D(n131),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][1]  (
	.SI(\regArr[10][0] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][1] ),
	.D(n130),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[10][0]  (
	.SI(\regArr[9][7] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[10][0] ),
	.D(n129),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][7]  (
	.SI(\regArr[6][6] ),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[6][7] ),
	.D(n104),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][6]  (
	.SI(\regArr[6][5] ),
	.SE(n234),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[6][6] ),
	.D(n103),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][5]  (
	.SI(\regArr[6][4] ),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[6][5] ),
	.D(n102),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][4]  (
	.SI(\regArr[6][3] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[6][4] ),
	.D(n101),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][3]  (
	.SI(\regArr[6][2] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[6][3] ),
	.D(n100),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][2]  (
	.SI(\regArr[6][1] ),
	.SE(n233),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[6][2] ),
	.D(n99),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][1]  (
	.SI(\regArr[6][0] ),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[6][1] ),
	.D(n98),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[6][0]  (
	.SI(\regArr[5][7] ),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[6][0] ),
	.D(n97),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][7]  (
	.SI(\regArr[12][6] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[12][7] ),
	.D(n152),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][6]  (
	.SI(\regArr[12][5] ),
	.SE(n234),
	.RN(RST),
	.Q(\regArr[12][6] ),
	.D(n151),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][5]  (
	.SI(\regArr[12][4] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[12][5] ),
	.D(n150),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][4]  (
	.SI(\regArr[12][3] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[12][4] ),
	.D(n149),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][3]  (
	.SI(\regArr[12][2] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[12][3] ),
	.D(n148),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][2]  (
	.SI(\regArr[12][1] ),
	.SE(n233),
	.RN(RST),
	.Q(\regArr[12][2] ),
	.D(n147),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][1]  (
	.SI(\regArr[12][0] ),
	.SE(n235),
	.RN(RST),
	.Q(\regArr[12][1] ),
	.D(n146),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[12][0]  (
	.SI(\regArr[11][7] ),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[12][0] ),
	.D(n145),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][7]  (
	.SI(\regArr[8][6] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][7] ),
	.D(n120),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][6]  (
	.SI(\regArr[8][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][6] ),
	.D(n119),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][5]  (
	.SI(\regArr[8][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][5] ),
	.D(n118),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][4]  (
	.SI(\regArr[8][3] ),
	.SE(n238),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][4] ),
	.D(n117),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][3]  (
	.SI(\regArr[8][2] ),
	.SE(n237),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][3] ),
	.D(n116),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][2]  (
	.SI(\regArr[8][1] ),
	.SE(n233),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][2] ),
	.D(n115),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][1]  (
	.SI(\regArr[8][0] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[8][1] ),
	.D(n114),
	.CK(REF_SCAN_CLK__L6_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[8][0]  (
	.SI(\regArr[7][7] ),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[8][0] ),
	.D(n113),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][7]  (
	.SI(\regArr[4][6] ),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[4][7] ),
	.D(n88),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][6]  (
	.SI(\regArr[4][5] ),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[4][6] ),
	.D(n87),
	.CK(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][5]  (
	.SI(\regArr[4][4] ),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(\regArr[4][5] ),
	.D(n86),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][4]  (
	.SI(\regArr[4][3] ),
	.SE(n238),
	.RN(RST),
	.Q(\regArr[4][4] ),
	.D(n85),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][3]  (
	.SI(\regArr[4][2] ),
	.SE(n237),
	.RN(RST),
	.Q(\regArr[4][3] ),
	.D(n84),
	.CK(REF_SCAN_CLK__L6_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][2]  (
	.SI(\regArr[4][1] ),
	.SE(n233),
	.RN(RST),
	.Q(\regArr[4][2] ),
	.D(n83),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][1]  (
	.SI(\regArr[4][0] ),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[4][1] ),
	.D(n82),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[4][0]  (
	.SI(REG3[7]),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(\regArr[4][0] ),
	.D(n81),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[7]  (
	.SI(RdData[6]),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[7]),
	.D(n47),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[6]  (
	.SI(RdData[5]),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[6]),
	.D(n46),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[5]  (
	.SI(RdData[4]),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[5]),
	.D(n45),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[4]  (
	.SI(RdData[3]),
	.SE(n233),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[4]),
	.D(n44),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[3]  (
	.SI(RdData[2]),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[3]),
	.D(n43),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[2]  (
	.SI(RdData[1]),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[2]),
	.D(n42),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[1]  (
	.SI(RdData[0]),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(RdData[1]),
	.D(n41),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[0]  (
	.SI(RdData_VLD),
	.SE(n234),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(RdData[0]),
	.D(n40),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RdData_VLD_reg (
	.SI(test_si1),
	.SE(n235),
	.RN(FE_OFN0_SYNC_SCAN_RST1),
	.Q(RdData_VLD),
	.D(n48),
	.CK(REF_SCAN_CLK__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][6]  (
	.SI(REG1[5]),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG1[6]),
	.D(n63),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][7]  (
	.SI(REG0[6]),
	.SE(n235),
	.RN(RST),
	.Q(REG0[7]),
	.D(n56),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][6]  (
	.SI(REG0[5]),
	.SE(n238),
	.RN(RST),
	.Q(REG0[6]),
	.D(n55),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][5]  (
	.SI(REG0[4]),
	.SE(n237),
	.RN(RST),
	.Q(REG0[5]),
	.D(n54),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][4]  (
	.SI(REG0[3]),
	.SE(n233),
	.RN(RST),
	.Q(REG0[4]),
	.D(n53),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][3]  (
	.SI(REG0[2]),
	.SE(n235),
	.RN(RST),
	.Q(REG0[3]),
	.D(n52),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][2]  (
	.SI(REG0[1]),
	.SE(n238),
	.RN(RST),
	.Q(REG0[2]),
	.D(n51),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][1]  (
	.SI(REG0[0]),
	.SE(n237),
	.RN(RST),
	.Q(REG0[1]),
	.D(n50),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[0][0]  (
	.SI(RdData[7]),
	.SE(n234),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG0[0]),
	.D(n49),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[2][1]  (
	.SI(REG2[0]),
	.SE(n234),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG2[1]),
	.D(n66),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \regArr_reg[2][0]  (
	.SN(FE_OFN1_SYNC_SCAN_RST1),
	.SI(REG1[7]),
	.SE(n235),
	.Q(REG2[0]),
	.D(n65),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][0]  (
	.SI(test_si2),
	.SE(n235),
	.RN(RST),
	.Q(REG3[0]),
	.D(n73),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][1]  (
	.SI(REG1[0]),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG1[1]),
	.D(n58),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][5]  (
	.SI(REG1[4]),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG1[5]),
	.D(n62),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][4]  (
	.SI(REG1[3]),
	.SE(n233),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG1[4]),
	.D(n61),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][7]  (
	.SI(REG1[6]),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG1[7]),
	.D(n64),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][3]  (
	.SI(REG1[2]),
	.SE(n235),
	.RN(RST),
	.Q(REG1[3]),
	.D(n60),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][2]  (
	.SI(REG1[1]),
	.SE(n238),
	.RN(RST),
	.Q(REG1[2]),
	.D(n59),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[1][0]  (
	.SI(REG0[7]),
	.SE(n234),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG1[0]),
	.D(n57),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \regArr_reg[3][5]  (
	.SN(RST),
	.SI(REG3[4]),
	.SE(n238),
	.Q(REG3[5]),
	.D(n78),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][7]  (
	.SI(REG3[6]),
	.SE(n237),
	.RN(RST),
	.Q(REG3[7]),
	.D(n80),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][6]  (
	.SI(REG3[5]),
	.SE(n234),
	.RN(RST),
	.Q(REG3[6]),
	.D(n79),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][3]  (
	.SI(REG3[2]),
	.SE(n238),
	.RN(RST),
	.Q(REG3[3]),
	.D(n76),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][2]  (
	.SI(REG3[1]),
	.SE(n237),
	.RN(RST),
	.Q(REG3[2]),
	.D(n75),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][4]  (
	.SI(REG3[3]),
	.SE(n235),
	.RN(RST),
	.Q(REG3[4]),
	.D(n77),
	.CK(REF_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[3][1]  (
	.SI(REG3[0]),
	.SE(n233),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG3[1]),
	.D(n74),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[2][4]  (
	.SI(REG2[3]),
	.SE(n235),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG2[4]),
	.D(n69),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[2][3]  (
	.SI(REG2[2]),
	.SE(n238),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG2[3]),
	.D(n68),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[2][6]  (
	.SI(REG2[5]),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG2[6]),
	.D(n71),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[2][2]  (
	.SI(REG2[1]),
	.SE(n237),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG2[2]),
	.D(n67),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regArr_reg[2][5]  (
	.SI(REG2[4]),
	.SE(n233),
	.RN(FE_OFN1_SYNC_SCAN_RST1),
	.Q(REG2[5]),
	.D(n70),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U239 (
	.Y(n236),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U240 (
	.Y(n233),
	.A(n236), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U241 (
	.Y(n234),
	.A(n236), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U242 (
	.Y(n235),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U243 (
	.Y(n237),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U244 (
	.Y(n238),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U245 (
	.Y(n239),
	.A(\regArr[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U246 (
	.Y(n240),
	.A(n239), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \regArr_reg[2][7]  (
	.SN(FE_OFN1_SYNC_SCAN_RST1),
	.SI(REG2[6]),
	.SE(n233),
	.Q(n242),
	.D(n72),
	.CK(REF_SCAN_CLK__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \regArr_reg[13][4]  (
	.SI(\regArr[13][3] ),
	.SE(n238),
	.RN(RST),
	.Q(FE_OFN6_SO_1_),
	.D(n157),
	.CK(REF_SCAN_CLK__L6_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U247 (
	.Y(n229),
	.A(n242), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U248 (
	.Y(REG2[7]),
	.A(n229), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPER_WIDTH8_test_1 (
	A, 
	B, 
	ALU_FUN, 
	ALU_CLK, 
	RST, 
	EN, 
	ALU_OUT, 
	OUT_VALID, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input ALU_CLK;
   input RST;
   input EN;
   output [15:0] ALU_OUT;
   output OUT_VALID;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN5_n35;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N132;
   wire N157;
   wire N158;
   wire N159;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire [15:0] ALU_OUT_Comb;

   // Module instantiations
   BUFX2M FE_OFC5_n35 (
	.Y(FE_OFN5_n35),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(n31),
	.B(n124),
	.AN(FE_OFN5_n35), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U7 (
	.Y(ALU_OUT_Comb[9]),
	.B0(n32),
	.A1N(n31),
	.A0N(N118), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U8 (
	.Y(ALU_OUT_Comb[10]),
	.B0(n32),
	.A1N(n31),
	.A0N(N119), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U9 (
	.Y(ALU_OUT_Comb[11]),
	.B0(n32),
	.A1N(n31),
	.A0N(N120), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U10 (
	.Y(ALU_OUT_Comb[12]),
	.B0(n32),
	.A1N(n31),
	.A0N(N121), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U11 (
	.Y(ALU_OUT_Comb[13]),
	.B0(n32),
	.A1N(n31),
	.A0N(N122), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U12 (
	.Y(ALU_OUT_Comb[14]),
	.B0(n32),
	.A1N(n31),
	.A0N(N123), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U13 (
	.Y(ALU_OUT_Comb[15]),
	.B0(n32),
	.A1N(n31),
	.A0N(N124), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U14 (
	.Y(n47),
	.B0(n101),
	.A1N(n105),
	.A0N(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U15 (
	.Y(n48),
	.B0(n101),
	.A1N(n99),
	.A0N(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U16 (
	.Y(n37),
	.B(n137),
	.AN(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U17 (
	.Y(n42),
	.B(n105),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(n50),
	.B(n105),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U20 (
	.Y(n41),
	.B(n137),
	.A(n107), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n137),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n138),
	.A(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n140),
	.A(n107), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U24 (
	.Y(n32),
	.B(n123),
	.A(EN), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n124),
	.A(EN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U26 (
	.Y(n49),
	.C(ALU_FUN[2]),
	.B(n139),
	.AN(n105), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U27 (
	.Y(n35),
	.C(n139),
	.B(ALU_FUN[2]),
	.A(n137), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U28 (
	.Y(n106),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U29 (
	.Y(n46),
	.C(ALU_FUN[3]),
	.B(n136),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U30 (
	.Y(n36),
	.C(ALU_FUN[3]),
	.B(n136),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U31 (
	.Y(n107),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n136),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(n105),
	.B(ALU_FUN[3]),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U34 (
	.Y(n100),
	.B(ALU_FUN[0]),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U35 (
	.Y(n91),
	.C(n99),
	.B(ALU_FUN[0]),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n139),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U37 (
	.Y(n101),
	.C(ALU_FUN[3]),
	.B(ALU_FUN[0]),
	.A(n106), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U38 (
	.Y(n99),
	.B(n139),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U39 (
	.Y(n90),
	.D(n136),
	.C(ALU_FUN[3]),
	.B(n99),
	.A(N159), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U40 (
	.Y(ALU_OUT_Comb[2]),
	.B0(n124),
	.A2(n77),
	.A1(n76),
	.A0(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U41 (
	.Y(n75),
	.B1(n37),
	.B0(N93),
	.A1(n50),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U42 (
	.Y(n77),
	.C0(n78),
	.B1(n133),
	.B0(n41),
	.A1(n138),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U43 (
	.Y(n76),
	.C1(n49),
	.C0(N127),
	.B1(n42),
	.B0(A[2]),
	.A1(FE_OFN5_n35),
	.A0(N111), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U44 (
	.Y(ALU_OUT_Comb[3]),
	.B0(n124),
	.A2(n71),
	.A1(n70),
	.A0(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U45 (
	.Y(n69),
	.B1(n37),
	.B0(N94),
	.A1(n50),
	.A0(N103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U46 (
	.Y(n71),
	.C0(n72),
	.B1(n132),
	.B0(n41),
	.A1(n138),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U47 (
	.Y(n70),
	.C1(n49),
	.C0(N128),
	.B1(n42),
	.B0(A[3]),
	.A1(FE_OFN5_n35),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U48 (
	.Y(ALU_OUT_Comb[4]),
	.B0(n124),
	.A2(n65),
	.A1(n64),
	.A0(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U49 (
	.Y(n63),
	.B1(n37),
	.B0(N95),
	.A1(n50),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U50 (
	.Y(n65),
	.C0(n66),
	.B1(n131),
	.B0(n41),
	.A1(A[5]),
	.A0(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U51 (
	.Y(n64),
	.C1(n49),
	.C0(N129),
	.B1(n42),
	.B0(A[4]),
	.A1(FE_OFN5_n35),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U52 (
	.Y(ALU_OUT_Comb[5]),
	.B0(n124),
	.A2(n59),
	.A1(n58),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U53 (
	.Y(n57),
	.B1(n37),
	.B0(N96),
	.A1(n50),
	.A0(N105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U54 (
	.Y(n59),
	.C0(n60),
	.B1(n130),
	.B0(n41),
	.A1(A[6]),
	.A0(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U55 (
	.Y(n58),
	.C1(n49),
	.C0(N130),
	.B1(n42),
	.B0(A[5]),
	.A1(FE_OFN5_n35),
	.A0(N114), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U56 (
	.Y(ALU_OUT_Comb[6]),
	.B0(n124),
	.A2(n53),
	.A1(n52),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U57 (
	.Y(n51),
	.B1(n37),
	.B0(N97),
	.A1(n50),
	.A0(N106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U58 (
	.Y(n53),
	.C0(n54),
	.B1(n129),
	.B0(n41),
	.A1(A[7]),
	.A0(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U59 (
	.Y(n52),
	.C1(n49),
	.C0(N131),
	.B1(A[6]),
	.B0(n42),
	.A1(FE_OFN5_n35),
	.A0(N115), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U60 (
	.Y(ALU_OUT_Comb[7]),
	.B0(n124),
	.A2(n40),
	.A1(n39),
	.A0(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U61 (
	.Y(n39),
	.B1(FE_OFN5_n35),
	.B0(N116),
	.A1(n49),
	.A0(N132), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U62 (
	.Y(n38),
	.B1(n37),
	.B0(N98),
	.A1(n50),
	.A0(N107), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U63 (
	.Y(n40),
	.C0(n43),
	.B1(A[7]),
	.B0(n42),
	.A1(n128),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U64 (
	.Y(ALU_OUT_Comb[0]),
	.B0(n124),
	.A2(n95),
	.A1(n94),
	.A0(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U65 (
	.Y(n93),
	.B1(n37),
	.B0(N91),
	.A1(n50),
	.A0(N100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U66 (
	.Y(n95),
	.C0(n97),
	.B0(n96),
	.A1(n135),
	.A0(n41), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U67 (
	.Y(n94),
	.C1(n49),
	.C0(N125),
	.B1(n42),
	.B0(A[0]),
	.A1(FE_OFN5_n35),
	.A0(N109), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U68 (
	.Y(ALU_OUT_Comb[1]),
	.B0(n124),
	.A2(n83),
	.A1(n82),
	.A0(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U69 (
	.Y(n83),
	.C0(n85),
	.B0(n84),
	.A1(n138),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U70 (
	.Y(n82),
	.C1(n42),
	.C0(A[1]),
	.B1(n134),
	.B0(n41),
	.A1(n49),
	.A0(N126), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U71 (
	.Y(n81),
	.C1(n50),
	.C0(N101),
	.B1(FE_OFN5_n35),
	.B0(N110),
	.A1(n37),
	.A0(N92), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U72 (
	.Y(ALU_OUT_Comb[8]),
	.B0(n124),
	.A1(n34),
	.A0(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U73 (
	.Y(n33),
	.B0(n123),
	.A1(n37),
	.A0(N99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U74 (
	.Y(n34),
	.B1(FE_OFN5_n35),
	.B0(N117),
	.A1N(n36),
	.A0N(n128), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U75 (
	.Y(n122),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U76 (
	.Y(n54),
	.C1(n130),
	.C0(n36),
	.B1(n56),
	.B0(B[6]),
	.A1(n122),
	.A0(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U77 (
	.Y(n56),
	.C0(n41),
	.B1(n129),
	.B0(n47),
	.A1(n46),
	.A0(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U78 (
	.Y(n55),
	.C0(n42),
	.B1(n48),
	.B0(A[6]),
	.A1(n129),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(n123),
	.A(n92), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U80 (
	.Y(n92),
	.C0(n47),
	.B0(n41),
	.A1(n50),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U82 (
	.Y(n134),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U83 (
	.Y(n135),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U84 (
	.Y(n129),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U85 (
	.Y(n128),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U86 (
	.Y(n132),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U87 (
	.Y(n133),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U88 (
	.Y(n130),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U89 (
	.Y(n131),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U90 (
	.Y(n78),
	.C1(n134),
	.C0(n36),
	.B1(n80),
	.B0(B[2]),
	.A1(n119),
	.A0(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U91 (
	.Y(n80),
	.C0(n41),
	.B1(n133),
	.B0(n47),
	.A1(n46),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U92 (
	.Y(n79),
	.C0(n42),
	.B1(n48),
	.B0(A[2]),
	.A1(n133),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U93 (
	.Y(n72),
	.C1(n133),
	.C0(n36),
	.B1(n74),
	.B0(B[3]),
	.A1(n121),
	.A0(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U94 (
	.Y(n74),
	.C0(n41),
	.B1(n132),
	.B0(n47),
	.A1(n46),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U95 (
	.Y(n73),
	.C0(n42),
	.B1(n48),
	.B0(A[3]),
	.A1(n132),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U96 (
	.Y(n66),
	.C1(n132),
	.C0(n36),
	.B1(n68),
	.B0(B[4]),
	.A1(n127),
	.A0(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n127),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U98 (
	.Y(n68),
	.C0(n41),
	.B1(n131),
	.B0(n47),
	.A1(n46),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U99 (
	.Y(n67),
	.C0(n42),
	.B1(n48),
	.B0(A[4]),
	.A1(n131),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U100 (
	.Y(n60),
	.C1(n131),
	.C0(n36),
	.B1(n62),
	.B0(B[5]),
	.A1(n126),
	.A0(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U101 (
	.Y(n126),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U102 (
	.Y(n62),
	.C0(n41),
	.B1(n130),
	.B0(n47),
	.A1(n46),
	.A0(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U103 (
	.Y(n61),
	.C0(n42),
	.B1(n48),
	.B0(A[5]),
	.A1(n130),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U104 (
	.Y(n43),
	.C1(n129),
	.C0(n36),
	.B1(n45),
	.B0(B[7]),
	.A1(n125),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U105 (
	.Y(n125),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U106 (
	.Y(n45),
	.C0(n41),
	.B1(n128),
	.B0(n47),
	.A1(A[7]),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U107 (
	.Y(n44),
	.C0(n42),
	.B1(n48),
	.B0(A[7]),
	.A1(n128),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n118),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U109 (
	.Y(n97),
	.B1(n134),
	.B0(n91),
	.A1N(B[0]),
	.A0(n98), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U110 (
	.Y(n98),
	.C0(n42),
	.B1(n48),
	.B0(A[0]),
	.A1(n135),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U111 (
	.Y(n85),
	.B1(n135),
	.B0(n36),
	.A1N(B[1]),
	.A0(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U112 (
	.Y(n86),
	.C0(n42),
	.B1(n48),
	.B0(A[1]),
	.A1(n134),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U113 (
	.Y(n120),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U114 (
	.Y(n96),
	.B0(n103),
	.A1(n102),
	.A0(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U115 (
	.Y(n103),
	.B0(n90),
	.A2(n104),
	.A1(ALU_FUN[3]),
	.A0(N157), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U116 (
	.Y(n102),
	.C0(n41),
	.B1(n135),
	.B0(n47),
	.A1(n46),
	.A0(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U117 (
	.Y(n104),
	.C(ALU_FUN[0]),
	.B(ALU_FUN[2]),
	.A(n139), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U118 (
	.Y(n84),
	.B0(n88),
	.A1(n87),
	.A0(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U119 (
	.Y(n88),
	.B0(n90),
	.A2(n89),
	.A1(ALU_FUN[3]),
	.A0(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U120 (
	.Y(n87),
	.C0(n41),
	.B1(n134),
	.B0(n47),
	.A1(n46),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U121 (
	.Y(n89),
	.C(n139),
	.B(ALU_FUN[2]),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U130 (
	.Y(n117),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U131 (
	.Y(n119),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U132 (
	.Y(n121),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U133 (
	.Y(n113),
	.B(B[7]),
	.A(n128), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U134 (
	.Y(n29),
	.B(A[4]),
	.AN(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U135 (
	.Y(n18),
	.B(B[4]),
	.AN(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U136 (
	.Y(n108),
	.B(n18),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U137 (
	.Y(n26),
	.B(A[3]),
	.A(n121), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U138 (
	.Y(n17),
	.B(A[2]),
	.A(n119), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U139 (
	.Y(n14),
	.B(A[0]),
	.A(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U140 (
	.Y(n28),
	.B(n119),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U141 (
	.Y(n23),
	.B(n28),
	.AN(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U142 (
	.Y(n15),
	.B0(B[1]),
	.A1(n134),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U143 (
	.Y(n16),
	.C0(n15),
	.B0(n23),
	.A1(n118),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U144 (
	.Y(n27),
	.B(n121),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U145 (
	.Y(n19),
	.B0(n27),
	.A2(n16),
	.A1(n17),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U146 (
	.Y(n111),
	.B(B[5]),
	.AN(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U147 (
	.Y(n20),
	.C0(n111),
	.B0(n18),
	.A1(n19),
	.A0(n108), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U148 (
	.Y(n30),
	.B(A[5]),
	.AN(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U149 (
	.Y(n110),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U150 (
	.Y(n21),
	.B1(n129),
	.B0(B[6]),
	.A2(n110),
	.A1(n30),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U151 (
	.Y(n114),
	.B(n128),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U152 (
	.Y(N159),
	.B0(n114),
	.A1(n21),
	.A0(n113), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U153 (
	.Y(n24),
	.B(n117),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U154 (
	.Y(n22),
	.B0(B[1]),
	.A1(n134),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U155 (
	.Y(n25),
	.C0(n22),
	.B0(n23),
	.A1(n134),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U156 (
	.Y(n109),
	.B0(n26),
	.A2(n27),
	.A1(n28),
	.A0(n120), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X1M U157 (
	.Y(n112),
	.C0(n29),
	.B0(n30),
	.A1N(n109),
	.A0(n108), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U158 (
	.Y(n115),
	.B1(n122),
	.B0(A[6]),
	.A2(n110),
	.A1(n111),
	.A0(n112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U159 (
	.Y(n116),
	.B0(n113),
	.A1N(n115),
	.A0(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U160 (
	.Y(N158),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U161 (
	.Y(N157),
	.B(N158),
	.A(N159), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[15]),
	.D(ALU_OUT_Comb[15]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[14]),
	.D(ALU_OUT_Comb[14]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[13]),
	.D(ALU_OUT_Comb[13]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[12]),
	.D(ALU_OUT_Comb[12]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[11]),
	.D(ALU_OUT_Comb[11]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[10]),
	.D(ALU_OUT_Comb[10]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[9]),
	.D(ALU_OUT_Comb[9]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[8]),
	.D(ALU_OUT_Comb[8]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[7]),
	.D(ALU_OUT_Comb[7]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[6]),
	.D(ALU_OUT_Comb[6]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[5]),
	.D(ALU_OUT_Comb[5]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[4]),
	.D(ALU_OUT_Comb[4]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[3]),
	.D(ALU_OUT_Comb[3]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[2]),
	.D(ALU_OUT_Comb[2]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[1]),
	.D(ALU_OUT_Comb[1]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[0]),
	.D(ALU_OUT_Comb[0]),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M OUT_VALID_reg (
	.SI(ALU_OUT[15]),
	.SE(test_se),
	.RN(RST),
	.Q(OUT_VALID),
	.D(EN),
	.CK(ALU_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPER_WIDTH8_DW_div_uns_0 div_47 (
	.a({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.b({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.quotient({ N132,
		N131,
		N130,
		N129,
		N128,
		N127,
		N126,
		N125 }),
	.n117(n117),
	.n119(n119),
	.n121(n121),
	.n125(n125),
	.n127(n127),
	.n126(n126),
	.n135(n135),
	.n134(n134),
	.n133(n133),
	.n132(n132),
	.n131(n131),
	.n130(n130),
	.n129(n129),
	.n122(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPER_WIDTH8_DW01_sub_0 sub_41 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.DIFF({ N108,
		N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101,
		N100 }),
	.n117(n117),
	.n119(n119),
	.n121(n121),
	.n125(n125),
	.n127(n127),
	.n126(n126),
	.n135(n135),
	.n122(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPER_WIDTH8_DW01_add_0 add_38 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.SUM({ N99,
		N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92,
		N91 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPER_WIDTH8_DW02_mult_0 mult_44 (
	.A({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.TC(1'b0),
	.PRODUCT({ N124,
		N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109 }),
	.n117(n117),
	.n119(n119),
	.n121(n121),
	.n125(n125),
	.n127(n127),
	.n126(n126),
	.n135(n135),
	.n134(n134),
	.n133(n133),
	.n132(n132),
	.n131(n131),
	.n130(n130),
	.n129(n129),
	.n128(n128),
	.n122(n122), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPER_WIDTH8_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n117, 
	n119, 
	n121, 
	n125, 
	n127, 
	n126, 
	n135, 
	n134, 
	n133, 
	n132, 
	n131, 
	n130, 
	n129, 
	n122, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n117;
   input n119;
   input n121;
   input n125;
   input n127;
   input n126;
   input n135;
   input n134;
   input n133;
   input n132;
   input n131;
   input n130;
   input n129;
   input n122;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[1][4] ;
   wire \u_div/CryTmp[1][5] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][4] ;
   wire \u_div/CryTmp[2][5] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[3][4] ;
   wire \u_div/CryTmp[3][5] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[4][4] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[6][2] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n5;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;

   // Module instantiations
   ADDFX2M \u_div/u_fa_PartRem_0_2_5  (
	.S(\u_div/SumTmp[2][5] ),
	.CO(\u_div/CryTmp[2][6] ),
	.CI(\u_div/CryTmp[2][5] ),
	.B(n13),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_3  (
	.S(\u_div/SumTmp[4][3] ),
	.CO(\u_div/CryTmp[4][4] ),
	.CI(\u_div/CryTmp[4][3] ),
	.B(n15),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_2  (
	.S(\u_div/SumTmp[5][2] ),
	.CO(\u_div/CryTmp[5][3] ),
	.CI(\u_div/CryTmp[5][2] ),
	.B(n16),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_6_1  (
	.S(\u_div/SumTmp[6][1] ),
	.CO(\u_div/CryTmp[6][2] ),
	.CI(\u_div/CryTmp[6][1] ),
	.B(n17),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_4  (
	.S(\u_div/SumTmp[3][4] ),
	.CO(\u_div/CryTmp[3][5] ),
	.CI(\u_div/CryTmp[3][4] ),
	.B(n14),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(n13),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(n12),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(n11),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/CryTmp[0][1] ),
	.B(n17),
	.A(\u_div/PartRem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_1  (
	.S(\u_div/SumTmp[1][1] ),
	.CO(\u_div/CryTmp[1][2] ),
	.CI(\u_div/CryTmp[1][1] ),
	.B(n17),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_1  (
	.S(\u_div/SumTmp[2][1] ),
	.CO(\u_div/CryTmp[2][2] ),
	.CI(\u_div/CryTmp[2][1] ),
	.B(n17),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_1  (
	.S(\u_div/SumTmp[3][1] ),
	.CO(\u_div/CryTmp[3][2] ),
	.CI(\u_div/CryTmp[3][1] ),
	.B(n17),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_1  (
	.S(\u_div/SumTmp[4][1] ),
	.CO(\u_div/CryTmp[4][2] ),
	.CI(\u_div/CryTmp[4][1] ),
	.B(n17),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_5_1  (
	.S(\u_div/SumTmp[5][1] ),
	.CO(\u_div/CryTmp[5][2] ),
	.CI(\u_div/CryTmp[5][1] ),
	.B(n17),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(n16),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(n15),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(n14),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_5  (
	.S(\u_div/SumTmp[1][5] ),
	.CO(\u_div/CryTmp[1][6] ),
	.CI(\u_div/CryTmp[1][5] ),
	.B(n13),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_4  (
	.S(\u_div/SumTmp[1][4] ),
	.CO(\u_div/CryTmp[1][5] ),
	.CI(\u_div/CryTmp[1][4] ),
	.B(n14),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_3  (
	.S(\u_div/SumTmp[1][3] ),
	.CO(\u_div/CryTmp[1][4] ),
	.CI(\u_div/CryTmp[1][3] ),
	.B(n15),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_4  (
	.S(\u_div/SumTmp[2][4] ),
	.CO(\u_div/CryTmp[2][5] ),
	.CI(\u_div/CryTmp[2][4] ),
	.B(n14),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_2  (
	.S(\u_div/SumTmp[1][2] ),
	.CO(\u_div/CryTmp[1][3] ),
	.CI(\u_div/CryTmp[1][2] ),
	.B(n16),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_3  (
	.S(\u_div/SumTmp[2][3] ),
	.CO(\u_div/CryTmp[2][4] ),
	.CI(\u_div/CryTmp[2][3] ),
	.B(n15),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_2_2  (
	.S(\u_div/SumTmp[2][2] ),
	.CO(\u_div/CryTmp[2][3] ),
	.CI(\u_div/CryTmp[2][2] ),
	.B(n16),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_3  (
	.S(\u_div/SumTmp[3][3] ),
	.CO(\u_div/CryTmp[3][4] ),
	.CI(\u_div/CryTmp[3][3] ),
	.B(n15),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_3_2  (
	.S(\u_div/SumTmp[3][2] ),
	.CO(\u_div/CryTmp[3][3] ),
	.CI(\u_div/CryTmp[3][2] ),
	.B(n16),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_4_2  (
	.S(\u_div/SumTmp[4][2] ),
	.CO(\u_div/CryTmp[4][3] ),
	.CI(\u_div/CryTmp[4][2] ),
	.B(n16),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M \u_div/u_fa_PartRem_0_1_6  (
	.S(\u_div/SumTmp[1][6] ),
	.CO(\u_div/CryTmp[1][7] ),
	.CI(\u_div/CryTmp[1][6] ),
	.B(n12),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(n18),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(\u_div/SumTmp[6][0] ),
	.B(a[6]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(\u_div/SumTmp[5][0] ),
	.B(a[5]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(\u_div/SumTmp[4][0] ),
	.B(a[4]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(\u_div/SumTmp[1][0] ),
	.B(a[1]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(\u_div/CryTmp[5][1] ),
	.B(n3),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n3),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n2),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U13 (
	.Y(\u_div/CryTmp[4][1] ),
	.B(n5),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n5),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(n7),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n7),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n8),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n8),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U21 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(n9),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n9),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(n10),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n10),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(n1),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n1),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n12),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n17),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n16),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n15),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n14),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n13),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n11),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U34 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][6] ),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U35 (
	.Y(\u_div/PartRem[2][6] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U36 (
	.Y(\u_div/PartRem[3][5] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U37 (
	.Y(\u_div/PartRem[4][4] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U38 (
	.Y(\u_div/PartRem[5][3] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U39 (
	.Y(\u_div/PartRem[6][2] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][1] ),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U40 (
	.Y(\u_div/PartRem[7][1] ),
	.S0(quotient[7]),
	.B(\u_div/SumTmp[7][0] ),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U41 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][5] ),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U42 (
	.Y(\u_div/PartRem[2][5] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U43 (
	.Y(\u_div/PartRem[3][4] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U44 (
	.Y(\u_div/PartRem[4][3] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][2] ),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U45 (
	.Y(\u_div/PartRem[5][2] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][1] ),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U46 (
	.Y(\u_div/PartRem[6][1] ),
	.S0(quotient[6]),
	.B(\u_div/SumTmp[6][0] ),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U47 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][4] ),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U48 (
	.Y(\u_div/PartRem[2][4] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U49 (
	.Y(\u_div/PartRem[3][3] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U50 (
	.Y(\u_div/PartRem[4][2] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][1] ),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U51 (
	.Y(\u_div/PartRem[5][1] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][0] ),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U52 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][3] ),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U53 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U54 (
	.Y(\u_div/PartRem[3][2] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][1] ),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U55 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][0] ),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U56 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][2] ),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U57 (
	.Y(\u_div/PartRem[2][2] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][1] ),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U58 (
	.Y(\u_div/PartRem[3][1] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][0] ),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U59 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][1] ),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U60 (
	.Y(\u_div/PartRem[2][1] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][0] ),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U61 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][0] ),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X1M U62 (
	.Y(quotient[7]),
	.D(n16),
	.C(n17),
	.B(n19),
	.A(\u_div/CryTmp[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U63 (
	.Y(quotient[6]),
	.C(\u_div/CryTmp[6][2] ),
	.B(n16),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U64 (
	.Y(quotient[5]),
	.B(n19),
	.A(\u_div/CryTmp[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U65 (
	.Y(n19),
	.B(n15),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U66 (
	.Y(quotient[4]),
	.B(n20),
	.A(\u_div/CryTmp[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U67 (
	.Y(n20),
	.C(n13),
	.B(n14),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X1M U68 (
	.Y(quotient[3]),
	.C(\u_div/CryTmp[3][5] ),
	.B(n13),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U69 (
	.Y(quotient[2]),
	.B(n21),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(n21),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U71 (
	.Y(quotient[1]),
	.B(n11),
	.A(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPER_WIDTH8_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n117, 
	n119, 
	n121, 
	n125, 
	n127, 
	n126, 
	n135, 
	n122, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n117;
   input n119;
   input n121;
   input n125;
   input n127;
   input n126;
   input n135;
   input n122;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n2),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n8),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n4),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n5),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n6),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n7),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n3),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U1 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(n3),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n9),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n7),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n6),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n5),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n4),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U8 (
	.Y(carry[1]),
	.B(n1),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n8),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n1),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n2),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U12 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPER_WIDTH8_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[0]),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPER_WIDTH8_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n117, 
	n119, 
	n121, 
	n125, 
	n127, 
	n126, 
	n135, 
	n134, 
	n133, 
	n132, 
	n131, 
	n130, 
	n129, 
	n128, 
	n122, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n117;
   input n119;
   input n121;
   input n125;
   input n127;
   input n126;
   input n135;
   input n134;
   input n133;
   input n132;
   input n131;
   input n130;
   input n129;
   input n128;
   input n122;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;

   // Module instantiations
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n8),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n9),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n7),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n6),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n5),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n4),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n3),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n22),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(PRODUCT[1]),
	.B(\ab[0][1] ),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n23),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n21),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n20),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n19),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n18),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U23 (
	.Y(\A1[6] ),
	.B(n17),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n17),
	.A(\SUMB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U25 (
	.Y(n11),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U26 (
	.Y(n12),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U27 (
	.Y(n13),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n14),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U30 (
	.Y(n16),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U31 (
	.Y(\SUMB[1][6] ),
	.B(n23),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(\SUMB[1][5] ),
	.B(n22),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U33 (
	.Y(\SUMB[1][4] ),
	.B(n21),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U34 (
	.Y(\SUMB[1][3] ),
	.B(n20),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][2] ),
	.B(n19),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U36 (
	.Y(\SUMB[1][1] ),
	.B(n18),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n32),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n33),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n38),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n39),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n36),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n37),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n34),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n35),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n25),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n31),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n29),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n28),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U49 (
	.Y(n24),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n27),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U51 (
	.Y(n26),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n30),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U54 (
	.Y(\ab[7][7] ),
	.B(n24),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][6] ),
	.B(n25),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][5] ),
	.B(n26),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][4] ),
	.B(n27),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][3] ),
	.B(n28),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][2] ),
	.B(n29),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][1] ),
	.B(n30),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[7][0] ),
	.B(n31),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[6][7] ),
	.B(n33),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][6] ),
	.B(n33),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][5] ),
	.B(n33),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][4] ),
	.B(n33),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][3] ),
	.B(n33),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][2] ),
	.B(n33),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][1] ),
	.B(n33),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][0] ),
	.B(n33),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[5][7] ),
	.B(n34),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][6] ),
	.B(n34),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][5] ),
	.B(n34),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][4] ),
	.B(n34),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][3] ),
	.B(n34),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][2] ),
	.B(n34),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][1] ),
	.B(n34),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][0] ),
	.B(n34),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[4][7] ),
	.B(n35),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][6] ),
	.B(n35),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][5] ),
	.B(n35),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][4] ),
	.B(n35),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][3] ),
	.B(n35),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][2] ),
	.B(n35),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][1] ),
	.B(n35),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][0] ),
	.B(n35),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[3][7] ),
	.B(n36),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][6] ),
	.B(n36),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][5] ),
	.B(n36),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][4] ),
	.B(n36),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][3] ),
	.B(n36),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][2] ),
	.B(n36),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][1] ),
	.B(n36),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][0] ),
	.B(n36),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[2][7] ),
	.B(n37),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][6] ),
	.B(n37),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][5] ),
	.B(n37),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][4] ),
	.B(n37),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][3] ),
	.B(n37),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][2] ),
	.B(n37),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][1] ),
	.B(n37),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][0] ),
	.B(n37),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[1][7] ),
	.B(n38),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][6] ),
	.B(n38),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][5] ),
	.B(n38),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][4] ),
	.B(n38),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][3] ),
	.B(n38),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][2] ),
	.B(n38),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][1] ),
	.B(n38),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][0] ),
	.B(n38),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[0][7] ),
	.B(n39),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][6] ),
	.B(n39),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][5] ),
	.B(n39),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][4] ),
	.B(n39),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][3] ),
	.B(n39),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][2] ),
	.B(n39),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(\ab[0][1] ),
	.B(n39),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U117 (
	.Y(PRODUCT[0]),
	.B(n39),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPER_WIDTH8_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n14,
		n16,
		n13,
		n15,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_OPER_WIDTH8_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   // Module instantiations
   AOI21BX2M U2 (
	.Y(n1),
	.B0N(n19),
	.A1(A[12]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(SUM[7]),
	.B(n8),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n8),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U6 (
	.Y(n15),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n9),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(SUM[6]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U9 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U10 (
	.Y(SUM[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U11 (
	.Y(SUM[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U12 (
	.Y(SUM[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U13 (
	.Y(SUM[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U14 (
	.Y(SUM[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U15 (
	.Y(SUM[9]),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(SUM[8]),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U18 (
	.Y(n14),
	.B(n17),
	.AN(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(n19),
	.B0(B[12]),
	.A1(n18),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U20 (
	.Y(SUM[12]),
	.C(n18),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U21 (
	.Y(n18),
	.B0N(n22),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U22 (
	.Y(SUM[11]),
	.B(n23),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U23 (
	.Y(n23),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(n20),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U25 (
	.Y(n22),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U26 (
	.Y(n21),
	.B0(n26),
	.A1(n25),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(SUM[10]),
	.B(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U28 (
	.Y(n25),
	.B0(n12),
	.A1N(n13),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U29 (
	.Y(n12),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(n13),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U31 (
	.Y(n10),
	.B0(n17),
	.A1(n16),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n17),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U33 (
	.Y(n16),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U34 (
	.Y(n27),
	.B(n26),
	.AN(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n26),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U36 (
	.Y(n24),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_GATE (
	CLK_EN, 
	CLK, 
	GATED_CLK, 
	VDD, 
	VSS);
   input CLK_EN;
   input CLK;
   output GATED_CLK;
   inout VDD;
   inout VSS;

   // Module instantiations
   TLATNCAX12M U0_TLATNCAX12M (
	.ECK(GATED_CLK),
	.E(CLK_EN),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_TOP (
	RST_N, 
	UART_CLK, 
	REF_CLK, 
	UART_RX_IN, 
	scan_clk, 
	scan_rst, 
	test_mode, 
	SE, 
	SI, 
	SO, 
	UART_TX_O, 
	parity_error, 
	framing_error, 
	VDD, 
	VSS);
   input RST_N;
   input UART_CLK;
   input REF_CLK;
   input UART_RX_IN;
   input scan_clk;
   input scan_rst;
   input test_mode;
   input SE;
   input [3:0] SI;
   output [3:0] SO;
   output UART_TX_O;
   output parity_error;
   output framing_error;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN22_SYNC_SCAN_RST2__Exclude_0_NET;
   wire FE_PHN21_SYNC_SCAN_RST2__Exclude_0_NET;
   wire FE_PHN20_SYNC_SCAN_RST2__Exclude_0_NET;
   wire FE_PHN19_SYNC_SCAN_RST2__Exclude_0_NET;
   wire FE_PHN18_SYNC_SCAN_RST2__Exclude_0_NET;
   wire FE_PHN17_SYNC_SCAN_RST2__Exclude_0_NET;
   wire FE_PHN14_SYNC_RST2__Exclude_0_NET;
   wire FE_PHN13_SYNC_RST2__Exclude_0_NET;
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L15_N0;
   wire scan_clk__L14_N0;
   wire scan_clk__L13_N1;
   wire scan_clk__L13_N0;
   wire scan_clk__L12_N1;
   wire scan_clk__L12_N0;
   wire scan_clk__L11_N1;
   wire scan_clk__L11_N0;
   wire scan_clk__L10_N1;
   wire scan_clk__L10_N0;
   wire scan_clk__L9_N1;
   wire scan_clk__L9_N0;
   wire scan_clk__L8_N1;
   wire scan_clk__L8_N0;
   wire scan_clk__L7_N1;
   wire scan_clk__L7_N0;
   wire scan_clk__L6_N1;
   wire scan_clk__L6_N0;
   wire scan_clk__L5_N1;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N1;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N1;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N2;
   wire scan_clk__L2_N1;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire REF_SCAN_CLK__L6_N13;
   wire REF_SCAN_CLK__L6_N12;
   wire REF_SCAN_CLK__L6_N11;
   wire REF_SCAN_CLK__L6_N10;
   wire REF_SCAN_CLK__L6_N9;
   wire REF_SCAN_CLK__L6_N8;
   wire REF_SCAN_CLK__L6_N7;
   wire REF_SCAN_CLK__L6_N6;
   wire REF_SCAN_CLK__L6_N5;
   wire REF_SCAN_CLK__L6_N4;
   wire REF_SCAN_CLK__L6_N3;
   wire REF_SCAN_CLK__L6_N2;
   wire REF_SCAN_CLK__L6_N1;
   wire REF_SCAN_CLK__L6_N0;
   wire REF_SCAN_CLK__L5_N13;
   wire REF_SCAN_CLK__L5_N12;
   wire REF_SCAN_CLK__L5_N11;
   wire REF_SCAN_CLK__L5_N10;
   wire REF_SCAN_CLK__L5_N9;
   wire REF_SCAN_CLK__L5_N8;
   wire REF_SCAN_CLK__L5_N7;
   wire REF_SCAN_CLK__L5_N6;
   wire REF_SCAN_CLK__L5_N5;
   wire REF_SCAN_CLK__L5_N4;
   wire REF_SCAN_CLK__L5_N3;
   wire REF_SCAN_CLK__L5_N2;
   wire REF_SCAN_CLK__L5_N1;
   wire REF_SCAN_CLK__L5_N0;
   wire REF_SCAN_CLK__L4_N4;
   wire REF_SCAN_CLK__L4_N3;
   wire REF_SCAN_CLK__L4_N2;
   wire REF_SCAN_CLK__L4_N1;
   wire REF_SCAN_CLK__L4_N0;
   wire REF_SCAN_CLK__L3_N1;
   wire REF_SCAN_CLK__L3_N0;
   wire REF_SCAN_CLK__L2_N1;
   wire REF_SCAN_CLK__L2_N0;
   wire REF_SCAN_CLK__L1_N0;
   wire CLK_ALU__L3_N0;
   wire CLK_ALU__L2_N0;
   wire CLK_ALU__L1_N0;
   wire UART_SCAN_CLK__L18_N1;
   wire UART_SCAN_CLK__L18_N0;
   wire UART_SCAN_CLK__L17_N0;
   wire UART_SCAN_CLK__L16_N0;
   wire UART_SCAN_CLK__L15_N0;
   wire UART_SCAN_CLK__L14_N0;
   wire UART_SCAN_CLK__L13_N2;
   wire UART_SCAN_CLK__L13_N1;
   wire UART_SCAN_CLK__L13_N0;
   wire UART_SCAN_CLK__L12_N1;
   wire UART_SCAN_CLK__L12_N0;
   wire UART_SCAN_CLK__L11_N1;
   wire UART_SCAN_CLK__L11_N0;
   wire UART_SCAN_CLK__L10_N1;
   wire UART_SCAN_CLK__L10_N0;
   wire UART_SCAN_CLK__L9_N3;
   wire UART_SCAN_CLK__L9_N2;
   wire UART_SCAN_CLK__L9_N1;
   wire UART_SCAN_CLK__L9_N0;
   wire UART_SCAN_CLK__L8_N2;
   wire UART_SCAN_CLK__L8_N1;
   wire UART_SCAN_CLK__L8_N0;
   wire UART_SCAN_CLK__L7_N2;
   wire UART_SCAN_CLK__L7_N1;
   wire UART_SCAN_CLK__L7_N0;
   wire UART_SCAN_CLK__L6_N1;
   wire UART_SCAN_CLK__L6_N0;
   wire UART_SCAN_CLK__L5_N0;
   wire UART_SCAN_CLK__L4_N0;
   wire UART_SCAN_CLK__L3_N1;
   wire UART_SCAN_CLK__L3_N0;
   wire UART_SCAN_CLK__L2_N0;
   wire UART_SCAN_CLK__L1_N0;
   wire SYNC_RST2__Exclude_0_NET;
   wire SYNC_SCAN_RST2__L1_N0;
   wire SYNC_SCAN_RST2__Exclude_0_NET;
   wire n20__L1_N0;
   wire n20__Exclude_0_NET;
   wire n21__Exclude_0_NET;
   wire RX_SCAN_CLK__L4_N1;
   wire RX_SCAN_CLK__L4_N0;
   wire RX_SCAN_CLK__L3_N0;
   wire RX_SCAN_CLK__L2_N0;
   wire RX_SCAN_CLK__L1_N0;
   wire TX_SCAN_CLK__L4_N1;
   wire TX_SCAN_CLK__L4_N0;
   wire TX_SCAN_CLK__L3_N0;
   wire TX_SCAN_CLK__L2_N0;
   wire TX_SCAN_CLK__L1_N0;
   wire FE_OFN8_SE;
   wire FE_OFN2_SYNC_SCAN_RST1;
   wire FE_OFN1_SYNC_SCAN_RST1;
   wire FE_OFN0_SYNC_SCAN_RST1;
   wire n36;
   wire REF_SCAN_CLK;
   wire UART_SCAN_CLK;
   wire RX_CLK;
   wire RX_SCAN_CLK;
   wire TX_CLK;
   wire TX_SCAN_CLK;
   wire RSTN_SCAN_RST;
   wire SYNC_RST1;
   wire SYNC_SCAN_RST1;
   wire SYNC_RST2;
   wire SYNC_SCAN_RST2;
   wire RX_VLD;
   wire RX_VLD_SYNC;
   wire WR_INC;
   wire RD_INC;
   wire FIFO_FULL;
   wire F_EMPTY;
   wire BUSY;
   wire ALU_OUT_VLD;
   wire RD_D_VLD;
   wire ALU_EN;
   wire GATE_EN;
   wire WrEn;
   wire RdEn;
   wire CLK_ALU;
   wire _1_net_;
   wire n2;
   wire n3;
   wire n4;
   wire n10;
   wire n11;
   wire n15;
   wire n16;
   wire n19;
   wire n20;
   wire n21;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire [7:0] RX_OUT_P;
   wire [7:0] RX_OUT_SYNC;
   wire [7:0] WR_DATA;
   wire [7:0] RD_DATA;
   wire [7:0] div_ratio;
   wire [7:0] UART_CONFIG;
   wire [7:0] Pre_div;
   wire [15:0] ALU_OUT;
   wire [7:0] Rd_D;
   wire [3:0] ALU_FUN;
   wire [3:0] Address;
   wire [7:0] Wr_D;
   wire [7:0] Op_A;
   wire [7:0] Op_B;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;
   wire SYNOPSYS_UNCONNECTED__3;

   assign SO[2] = UART_CONFIG[7] ;

   // Module instantiations
   CLKBUFX8M FE_PHC22_SYNC_SCAN_RST2__Exclude_0_NET (
	.Y(FE_PHN21_SYNC_SCAN_RST2__Exclude_0_NET),
	.A(FE_PHN22_SYNC_SCAN_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_PHC21_SYNC_SCAN_RST2__Exclude_0_NET (
	.Y(FE_PHN20_SYNC_SCAN_RST2__Exclude_0_NET),
	.A(FE_PHN21_SYNC_SCAN_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_PHC20_SYNC_SCAN_RST2__Exclude_0_NET (
	.Y(FE_PHN19_SYNC_SCAN_RST2__Exclude_0_NET),
	.A(FE_PHN20_SYNC_SCAN_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_PHC19_SYNC_SCAN_RST2__Exclude_0_NET (
	.Y(FE_PHN18_SYNC_SCAN_RST2__Exclude_0_NET),
	.A(FE_PHN19_SYNC_SCAN_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_PHC18_SYNC_SCAN_RST2__Exclude_0_NET (
	.Y(FE_PHN17_SYNC_SCAN_RST2__Exclude_0_NET),
	.A(FE_PHN18_SYNC_SCAN_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_PHC17_SYNC_SCAN_RST2__Exclude_0_NET (
	.Y(SYNC_SCAN_RST2__Exclude_0_NET),
	.A(FE_PHN17_SYNC_SCAN_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC14_SYNC_RST2__Exclude_0_NET (
	.Y(FE_PHN13_SYNC_RST2__Exclude_0_NET),
	.A(FE_PHN14_SYNC_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC13_SYNC_RST2__Exclude_0_NET (
	.Y(SYNC_RST2__Exclude_0_NET),
	.A(FE_PHN13_SYNC_RST2__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M REF_CLK__L2_I0 (
	.Y(REF_CLK__L2_N0),
	.A(REF_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M REF_CLK__L1_I0 (
	.Y(REF_CLK__L1_N0),
	.A(REF_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_CLK__L2_I0 (
	.Y(UART_CLK__L2_N0),
	.A(UART_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_CLK__L1_I0 (
	.Y(UART_CLK__L1_N0),
	.A(UART_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M scan_clk__L15_I0 (
	.Y(scan_clk__L15_N0),
	.A(scan_clk__L14_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L14_I0 (
	.Y(scan_clk__L14_N0),
	.A(scan_clk__L13_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L13_I1 (
	.Y(scan_clk__L13_N1),
	.A(scan_clk__L12_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M scan_clk__L13_I0 (
	.Y(scan_clk__L13_N0),
	.A(scan_clk__L12_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L12_I1 (
	.Y(scan_clk__L12_N1),
	.A(scan_clk__L11_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L12_I0 (
	.Y(scan_clk__L12_N0),
	.A(scan_clk__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L11_I1 (
	.Y(scan_clk__L11_N1),
	.A(scan_clk__L10_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L11_I0 (
	.Y(scan_clk__L11_N0),
	.A(scan_clk__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L10_I1 (
	.Y(scan_clk__L10_N1),
	.A(scan_clk__L9_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L10_I0 (
	.Y(scan_clk__L10_N0),
	.A(scan_clk__L9_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L9_I1 (
	.Y(scan_clk__L9_N1),
	.A(scan_clk__L8_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L9_I0 (
	.Y(scan_clk__L9_N0),
	.A(scan_clk__L8_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L8_I1 (
	.Y(scan_clk__L8_N1),
	.A(scan_clk__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L8_I0 (
	.Y(scan_clk__L8_N0),
	.A(scan_clk__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L7_I1 (
	.Y(scan_clk__L7_N1),
	.A(scan_clk__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L7_I0 (
	.Y(scan_clk__L7_N0),
	.A(scan_clk__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L6_I1 (
	.Y(scan_clk__L6_N1),
	.A(scan_clk__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L6_I0 (
	.Y(scan_clk__L6_N0),
	.A(scan_clk__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L5_I1 (
	.Y(scan_clk__L5_N1),
	.A(scan_clk__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L5_I0 (
	.Y(scan_clk__L5_N0),
	.A(scan_clk__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L4_I1 (
	.Y(scan_clk__L4_N1),
	.A(scan_clk__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L4_I0 (
	.Y(scan_clk__L4_N0),
	.A(scan_clk__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L3_I1 (
	.Y(scan_clk__L3_N1),
	.A(scan_clk__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L3_I0 (
	.Y(scan_clk__L3_N0),
	.A(scan_clk__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M scan_clk__L2_I2 (
	.Y(scan_clk__L2_N2),
	.A(scan_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX32M scan_clk__L2_I1 (
	.Y(scan_clk__L2_N1),
	.A(scan_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M scan_clk__L2_I0 (
	.Y(scan_clk__L2_N0),
	.A(scan_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk__L1_I0 (
	.Y(scan_clk__L1_N0),
	.A(scan_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I13 (
	.Y(REF_SCAN_CLK__L6_N13),
	.A(REF_SCAN_CLK__L5_N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I12 (
	.Y(REF_SCAN_CLK__L6_N12),
	.A(REF_SCAN_CLK__L5_N12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I11 (
	.Y(REF_SCAN_CLK__L6_N11),
	.A(REF_SCAN_CLK__L5_N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I10 (
	.Y(REF_SCAN_CLK__L6_N10),
	.A(REF_SCAN_CLK__L5_N10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I9 (
	.Y(REF_SCAN_CLK__L6_N9),
	.A(REF_SCAN_CLK__L5_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I8 (
	.Y(REF_SCAN_CLK__L6_N8),
	.A(REF_SCAN_CLK__L5_N8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I7 (
	.Y(REF_SCAN_CLK__L6_N7),
	.A(REF_SCAN_CLK__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I6 (
	.Y(REF_SCAN_CLK__L6_N6),
	.A(REF_SCAN_CLK__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I5 (
	.Y(REF_SCAN_CLK__L6_N5),
	.A(REF_SCAN_CLK__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I4 (
	.Y(REF_SCAN_CLK__L6_N4),
	.A(REF_SCAN_CLK__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I3 (
	.Y(REF_SCAN_CLK__L6_N3),
	.A(REF_SCAN_CLK__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I2 (
	.Y(REF_SCAN_CLK__L6_N2),
	.A(REF_SCAN_CLK__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I1 (
	.Y(REF_SCAN_CLK__L6_N1),
	.A(REF_SCAN_CLK__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L6_I0 (
	.Y(REF_SCAN_CLK__L6_N0),
	.A(REF_SCAN_CLK__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I13 (
	.Y(REF_SCAN_CLK__L5_N13),
	.A(REF_SCAN_CLK__L4_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I12 (
	.Y(REF_SCAN_CLK__L5_N12),
	.A(REF_SCAN_CLK__L4_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I11 (
	.Y(REF_SCAN_CLK__L5_N11),
	.A(REF_SCAN_CLK__L4_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I10 (
	.Y(REF_SCAN_CLK__L5_N10),
	.A(REF_SCAN_CLK__L4_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I9 (
	.Y(REF_SCAN_CLK__L5_N9),
	.A(REF_SCAN_CLK__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I8 (
	.Y(REF_SCAN_CLK__L5_N8),
	.A(REF_SCAN_CLK__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I7 (
	.Y(REF_SCAN_CLK__L5_N7),
	.A(REF_SCAN_CLK__L4_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I6 (
	.Y(REF_SCAN_CLK__L5_N6),
	.A(REF_SCAN_CLK__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I5 (
	.Y(REF_SCAN_CLK__L5_N5),
	.A(REF_SCAN_CLK__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I4 (
	.Y(REF_SCAN_CLK__L5_N4),
	.A(REF_SCAN_CLK__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I3 (
	.Y(REF_SCAN_CLK__L5_N3),
	.A(REF_SCAN_CLK__L4_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I2 (
	.Y(REF_SCAN_CLK__L5_N2),
	.A(REF_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I1 (
	.Y(REF_SCAN_CLK__L5_N1),
	.A(REF_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L5_I0 (
	.Y(REF_SCAN_CLK__L5_N0),
	.A(REF_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L4_I4 (
	.Y(REF_SCAN_CLK__L4_N4),
	.A(REF_SCAN_CLK__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L4_I3 (
	.Y(REF_SCAN_CLK__L4_N3),
	.A(REF_SCAN_CLK__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L4_I2 (
	.Y(REF_SCAN_CLK__L4_N2),
	.A(REF_SCAN_CLK__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L4_I1 (
	.Y(REF_SCAN_CLK__L4_N1),
	.A(REF_SCAN_CLK__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L4_I0 (
	.Y(REF_SCAN_CLK__L4_N0),
	.A(REF_SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M REF_SCAN_CLK__L3_I1 (
	.Y(REF_SCAN_CLK__L3_N1),
	.A(REF_SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX24M REF_SCAN_CLK__L3_I0 (
	.Y(REF_SCAN_CLK__L3_N0),
	.A(REF_SCAN_CLK__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX14M REF_SCAN_CLK__L2_I1 (
	.Y(REF_SCAN_CLK__L2_N1),
	.A(REF_SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M REF_SCAN_CLK__L2_I0 (
	.Y(REF_SCAN_CLK__L2_N0),
	.A(REF_SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M REF_SCAN_CLK__L1_I0 (
	.Y(REF_SCAN_CLK__L1_N0),
	.A(REF_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M CLK_ALU__L3_I0 (
	.Y(CLK_ALU__L3_N0),
	.A(CLK_ALU__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M CLK_ALU__L2_I0 (
	.Y(CLK_ALU__L2_N0),
	.A(CLK_ALU__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M CLK_ALU__L1_I0 (
	.Y(CLK_ALU__L1_N0),
	.A(CLK_ALU), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L18_I1 (
	.Y(UART_SCAN_CLK__L18_N1),
	.A(UART_SCAN_CLK__L17_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L18_I0 (
	.Y(UART_SCAN_CLK__L18_N0),
	.A(UART_SCAN_CLK__L17_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_SCAN_CLK__L17_I0 (
	.Y(UART_SCAN_CLK__L17_N0),
	.A(UART_SCAN_CLK__L16_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_SCAN_CLK__L16_I0 (
	.Y(UART_SCAN_CLK__L16_N0),
	.A(UART_SCAN_CLK__L15_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M UART_SCAN_CLK__L15_I0 (
	.Y(UART_SCAN_CLK__L15_N0),
	.A(UART_SCAN_CLK__L14_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L14_I0 (
	.Y(UART_SCAN_CLK__L14_N0),
	.A(UART_SCAN_CLK__L13_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L13_I2 (
	.Y(UART_SCAN_CLK__L13_N2),
	.A(UART_SCAN_CLK__L12_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L13_I1 (
	.Y(UART_SCAN_CLK__L13_N1),
	.A(UART_SCAN_CLK__L12_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L13_I0 (
	.Y(UART_SCAN_CLK__L13_N0),
	.A(UART_SCAN_CLK__L12_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L12_I1 (
	.Y(UART_SCAN_CLK__L12_N1),
	.A(UART_SCAN_CLK__L11_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M UART_SCAN_CLK__L12_I0 (
	.Y(UART_SCAN_CLK__L12_N0),
	.A(UART_SCAN_CLK__L11_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L11_I1 (
	.Y(UART_SCAN_CLK__L11_N1),
	.A(UART_SCAN_CLK__L10_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_SCAN_CLK__L11_I0 (
	.Y(UART_SCAN_CLK__L11_N0),
	.A(UART_SCAN_CLK__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L10_I1 (
	.Y(UART_SCAN_CLK__L10_N1),
	.A(UART_SCAN_CLK__L9_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M UART_SCAN_CLK__L10_I0 (
	.Y(UART_SCAN_CLK__L10_N0),
	.A(UART_SCAN_CLK__L9_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L9_I3 (
	.Y(UART_SCAN_CLK__L9_N3),
	.A(UART_SCAN_CLK__L8_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L9_I2 (
	.Y(UART_SCAN_CLK__L9_N2),
	.A(UART_SCAN_CLK__L8_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L9_I1 (
	.Y(UART_SCAN_CLK__L9_N1),
	.A(UART_SCAN_CLK__L8_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M UART_SCAN_CLK__L9_I0 (
	.Y(UART_SCAN_CLK__L9_N0),
	.A(UART_SCAN_CLK__L8_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_SCAN_CLK__L8_I2 (
	.Y(UART_SCAN_CLK__L8_N2),
	.A(UART_SCAN_CLK__L7_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L8_I1 (
	.Y(UART_SCAN_CLK__L8_N1),
	.A(UART_SCAN_CLK__L7_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L8_I0 (
	.Y(UART_SCAN_CLK__L8_N0),
	.A(UART_SCAN_CLK__L7_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M UART_SCAN_CLK__L7_I2 (
	.Y(UART_SCAN_CLK__L7_N2),
	.A(UART_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L7_I1 (
	.Y(UART_SCAN_CLK__L7_N1),
	.A(UART_SCAN_CLK__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L7_I0 (
	.Y(UART_SCAN_CLK__L7_N0),
	.A(UART_SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L6_I1 (
	.Y(UART_SCAN_CLK__L6_N1),
	.A(UART_SCAN_CLK__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M UART_SCAN_CLK__L6_I0 (
	.Y(UART_SCAN_CLK__L6_N0),
	.A(UART_SCAN_CLK__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L5_I0 (
	.Y(UART_SCAN_CLK__L5_N0),
	.A(UART_SCAN_CLK__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L4_I0 (
	.Y(UART_SCAN_CLK__L4_N0),
	.A(UART_SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX16M UART_SCAN_CLK__L3_I1 (
	.Y(UART_SCAN_CLK__L3_N1),
	.A(UART_SCAN_CLK__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX20M UART_SCAN_CLK__L3_I0 (
	.Y(UART_SCAN_CLK__L3_N0),
	.A(UART_SCAN_CLK__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX24M UART_SCAN_CLK__L2_I0 (
	.Y(UART_SCAN_CLK__L2_N0),
	.A(UART_SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M UART_SCAN_CLK__L1_I0 (
	.Y(UART_SCAN_CLK__L1_N0),
	.A(UART_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M SYNC_RST2__Exclude_0 (
	.Y(FE_PHN14_SYNC_RST2__Exclude_0_NET),
	.A(SYNC_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M SYNC_SCAN_RST2__L1_I0 (
	.Y(SYNC_SCAN_RST2__L1_N0),
	.A(SYNC_SCAN_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M SYNC_SCAN_RST2__Exclude_0 (
	.Y(FE_PHN22_SYNC_SCAN_RST2__Exclude_0_NET),
	.A(SYNC_SCAN_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M n20__L1_I0 (
	.Y(n20__L1_N0),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M n20__Exclude_0 (
	.Y(n20__Exclude_0_NET),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M n21__Exclude_0 (
	.Y(n21__Exclude_0_NET),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M RX_SCAN_CLK__L4_I1 (
	.Y(RX_SCAN_CLK__L4_N1),
	.A(RX_SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M RX_SCAN_CLK__L4_I0 (
	.Y(RX_SCAN_CLK__L4_N0),
	.A(RX_SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M RX_SCAN_CLK__L3_I0 (
	.Y(RX_SCAN_CLK__L3_N0),
	.A(RX_SCAN_CLK__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M RX_SCAN_CLK__L2_I0 (
	.Y(RX_SCAN_CLK__L2_N0),
	.A(RX_SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M RX_SCAN_CLK__L1_I0 (
	.Y(RX_SCAN_CLK__L1_N0),
	.A(RX_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M TX_SCAN_CLK__L4_I1 (
	.Y(TX_SCAN_CLK__L4_N1),
	.A(TX_SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M TX_SCAN_CLK__L4_I0 (
	.Y(TX_SCAN_CLK__L4_N0),
	.A(TX_SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M TX_SCAN_CLK__L3_I0 (
	.Y(TX_SCAN_CLK__L3_N0),
	.A(TX_SCAN_CLK__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M TX_SCAN_CLK__L2_I0 (
	.Y(TX_SCAN_CLK__L2_N0),
	.A(TX_SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX12M TX_SCAN_CLK__L1_I0 (
	.Y(TX_SCAN_CLK__L1_N0),
	.A(TX_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC8_SE (
	.Y(FE_OFN8_SE),
	.A(SE), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC2_SYNC_SCAN_RST1 (
	.Y(FE_OFN2_SYNC_SCAN_RST1),
	.A(FE_OFN0_SYNC_SCAN_RST1), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC1_SYNC_SCAN_RST1 (
	.Y(FE_OFN1_SYNC_SCAN_RST1),
	.A(FE_OFN0_SYNC_SCAN_RST1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC0_SYNC_SCAN_RST1 (
	.Y(FE_OFN0_SYNC_SCAN_RST1),
	.A(SYNC_SCAN_RST1), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U4 (
	.Y(n3),
	.A(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U5 (
	.Y(n4),
	.A(Address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U7 (
	.Y(_1_net_),
	.B(n2),
	.A(GATE_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U11 (
	.Y(n2),
	.A(test_mode), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U19 (
	.Y(n25),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n26),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U21 (
	.Y(n27),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U22 (
	.Y(n28),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U23 (
	.Y(n29),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U24 (
	.Y(n30),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U25 (
	.Y(n31),
	.A(SE), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U26 (
	.Y(n32),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U27 (
	.Y(n33),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U28 (
	.Y(n34),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U29 (
	.Y(n35),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_1 U0_mux2X1 (
	.IN_0(REF_CLK__L2_N0),
	.IN_1(scan_clk__L13_N0),
	.SEL(n2),
	.OUT(REF_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_4 U1_mux2X1 (
	.IN_0(UART_CLK__L2_N0),
	.IN_1(scan_clk__L2_N0),
	.SEL(n2),
	.OUT(UART_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_3 U2_mux2X1 (
	.IN_0(RX_CLK),
	.IN_1(scan_clk__L15_N0),
	.SEL(n2),
	.OUT(RX_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_2 U3_mux2X1 (
	.IN_0(TX_CLK),
	.IN_1(scan_clk__L15_N0),
	.SEL(n2),
	.OUT(TX_SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_0 U4_mux2X1 (
	.IN_0(RST_N),
	.IN_1(scan_rst),
	.SEL(n2),
	.OUT(RSTN_SCAN_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_6 U5_mux2X1 (
	.IN_0(SYNC_RST1),
	.IN_1(scan_rst),
	.SEL(n2),
	.OUT(SYNC_SCAN_RST1), 
	.VDD(VDD), 
	.VSS(VSS));
   mux2X1_5 U6_mux2X1 (
	.IN_0(SYNC_RST2),
	.IN_1(scan_rst),
	.SEL(n2),
	.OUT(SYNC_SCAN_RST2), 
	.VDD(VDD), 
	.VSS(VSS));
   RST_SYNC_test_0 RST_SYNC1_INST (
	.CLK(REF_SCAN_CLK__L6_N0),
	.RST(RSTN_SCAN_RST),
	.SYNC_RST(SYNC_RST1),
	.test_si(n11),
	.test_se(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   RST_SYNC_test_1 RST_SYNC2_INST (
	.CLK(UART_SCAN_CLK__L18_N0),
	.RST(RSTN_SCAN_RST),
	.SYNC_RST(SYNC_RST2),
	.test_si(SYNC_RST1),
	.test_se(n28),
	.UART_SCAN_CLK__L3_N1(UART_SCAN_CLK__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   DataSynchronizer_BUS_WIDTH8_test_1 DATA_SYNC_INST (
	.Unsync_bus({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.bus_enable(RX_VLD),
	.CLK(REF_SCAN_CLK__L6_N5),
	.RST(FE_OFN1_SYNC_SCAN_RST1),
	.sync_bus({ RX_OUT_SYNC[7],
		RX_OUT_SYNC[6],
		RX_OUT_SYNC[5],
		RX_OUT_SYNC[4],
		RX_OUT_SYNC[3],
		RX_OUT_SYNC[2],
		RX_OUT_SYNC[1],
		RX_OUT_SYNC[0] }),
	.enable_pulse(RX_VLD_SYNC),
	.test_si(n20__Exclude_0_NET),
	.test_so(n19),
	.test_se(n28),
	.FE_OFN2_SYNC_SCAN_RST1(FE_OFN2_SYNC_SCAN_RST1), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_TOP_DATA_WIDTH8_test_1 FIFO_INST (
	.wclk(REF_SCAN_CLK__L6_N10),
	.rclk(TX_SCAN_CLK__L4_N0),
	.wrst_n(FE_OFN0_SYNC_SCAN_RST1),
	.rrst_n(SYNC_SCAN_RST2__Exclude_0_NET),
	.winc(WR_INC),
	.rinc(RD_INC),
	.wdata({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.rdata({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.wfull(FIFO_FULL),
	.empty(F_EMPTY),
	.test_si2(SI[2]),
	.test_si1(n19),
	.test_so2(n16),
	.test_so1(SO[3]),
	.test_se(FE_OFN8_SE),
	.FE_OFN2_SYNC_SCAN_RST1(FE_OFN2_SYNC_SCAN_RST1),
	.REF_SCAN_CLK__L6_N11(REF_SCAN_CLK__L6_N11),
	.REF_SCAN_CLK__L6_N12(REF_SCAN_CLK__L6_N12),
	.REF_SCAN_CLK__L6_N13(REF_SCAN_CLK__L6_N13),
	.REF_SCAN_CLK__L6_N4(REF_SCAN_CLK__L6_N4),
	.REF_SCAN_CLK__L6_N5(REF_SCAN_CLK__L6_N5),
	.REF_SCAN_CLK__L6_N6(REF_SCAN_CLK__L6_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   PULSE_GEN_test_1 PLSE_GEN_INST (
	.clk(TX_SCAN_CLK__L4_N0),
	.rst(SYNC_SCAN_RST2__Exclude_0_NET),
	.lvl_sig(BUSY),
	.pulse_sig(RD_INC),
	.test_si(n16),
	.test_so(n15),
	.test_se(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_test_1 CLK_DIV_TX_INST (
	.i_ref_clk(UART_SCAN_CLK__L13_N1),
	.i_rst_n(SYNC_SCAN_RST2__Exclude_0_NET),
	.i_clk_en(1'b1),
	.i_div_ratio({ div_ratio[7],
		div_ratio[6],
		div_ratio[5],
		div_ratio[4],
		div_ratio[3],
		div_ratio[2],
		div_ratio[1],
		div_ratio[0] }),
	.o_div_clk(TX_CLK),
	.test_si(n21__Exclude_0_NET),
	.test_so(n20),
	.test_se(n35),
	.n20__Exclude_0_NET(n20__Exclude_0_NET),
	.n20__L1_N0(n20__L1_N0),
	.SYNC_SCAN_RST2__L1_N0(SYNC_SCAN_RST2__L1_N0),
	.UART_SCAN_CLK__L18_N0(UART_SCAN_CLK__L18_N0),
	.UART_SCAN_CLK__L9_N3(UART_SCAN_CLK__L9_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKDIV_MUX PRE_MUX_INST (
	.IN({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2] }),
	.OUT({ SYNOPSYS_UNCONNECTED__0,
		SYNOPSYS_UNCONNECTED__1,
		SYNOPSYS_UNCONNECTED__2,
		SYNOPSYS_UNCONNECTED__3,
		Pre_div[3],
		Pre_div[2],
		Pre_div[1],
		Pre_div[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
   ClkDiv_test_0 CLK_DIV_RX_INST (
	.i_ref_clk(UART_SCAN_CLK__L13_N0),
	.i_rst_n(SYNC_SCAN_RST2__L1_N0),
	.i_clk_en(1'b1),
	.i_div_ratio({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		Pre_div[3],
		Pre_div[2],
		Pre_div[1],
		Pre_div[0] }),
	.o_div_clk(RX_CLK),
	.test_si(ALU_OUT_VLD),
	.test_so(n21),
	.test_se(n26),
	.n21__Exclude_0_NET(n21__Exclude_0_NET),
	.UART_SCAN_CLK__L18_N1(UART_SCAN_CLK__L18_N1),
	.UART_SCAN_CLK__L9_N2(UART_SCAN_CLK__L9_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_DATA_WIDTH8_test_1 UART_INST (
	.RST(SYNC_SCAN_RST2__Exclude_0_NET),
	.TX_CLK(TX_SCAN_CLK__L4_N0),
	.RX_CLK(RX_SCAN_CLK__L4_N0),
	.RX_IN_S(UART_RX_IN),
	.RX_OUT_P({ RX_OUT_P[7],
		RX_OUT_P[6],
		RX_OUT_P[5],
		RX_OUT_P[4],
		RX_OUT_P[3],
		RX_OUT_P[2],
		RX_OUT_P[1],
		RX_OUT_P[0] }),
	.RX_OUT_V(RX_VLD),
	.TX_IN_P({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }),
	.TX_IN_V(F_EMPTY),
	.TX_OUT_S(n36),
	.TX_OUT_V(BUSY),
	.Prescale({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2] }),
	.parity_enable(UART_CONFIG[0]),
	.parity_type(UART_CONFIG[1]),
	.parity_error(parity_error),
	.framing_error(framing_error),
	.test_si(n10),
	.test_se(FE_OFN8_SE),
	.TX_SCAN_CLK__L4_N1(TX_SCAN_CLK__L4_N1),
	.RX_SCAN_CLK__L4_N1(RX_SCAN_CLK__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SYS_CTRL_test_1 SYS_CTRL_INST (
	.clk(REF_SCAN_CLK__L6_N3),
	.rst_n(FE_OFN0_SYNC_SCAN_RST1),
	.RX_P_Data({ RX_OUT_SYNC[7],
		RX_OUT_SYNC[6],
		RX_OUT_SYNC[5],
		RX_OUT_SYNC[4],
		RX_OUT_SYNC[3],
		RX_OUT_SYNC[2],
		RX_OUT_SYNC[1],
		RX_OUT_SYNC[0] }),
	.RX_D_VLD(RX_VLD_SYNC),
	.RdData({ Rd_D[7],
		Rd_D[6],
		Rd_D[5],
		Rd_D[4],
		Rd_D[3],
		Rd_D[2],
		Rd_D[1],
		Rd_D[0] }),
	.RdData_Valid(RD_D_VLD),
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }),
	.OUT_Valid(ALU_OUT_VLD),
	.FIFO_FULL(FIFO_FULL),
	.Address({ Address[3],
		Address[2],
		Address[1],
		Address[0] }),
	.WrEn(WrEn),
	.RdEn(RdEn),
	.WrData({ Wr_D[7],
		Wr_D[6],
		Wr_D[5],
		Wr_D[4],
		Wr_D[3],
		Wr_D[2],
		Wr_D[1],
		Wr_D[0] }),
	.ALU_EN(ALU_EN),
	.ALU_FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }),
	.CLK_EN(GATE_EN),
	.WR_DATA({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }),
	.WR_INC(WR_INC),
	.test_si(SYNC_RST2__Exclude_0_NET),
	.test_so(n10),
	.test_se(n34),
	.FE_OFN2_SYNC_SCAN_RST1(FE_OFN2_SYNC_SCAN_RST1),
	.REF_SCAN_CLK__L6_N4(REF_SCAN_CLK__L6_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   RegFile_WIDTH8_DEPTH16_test_1 REG_FILE_INST (
	.CLK(REF_SCAN_CLK__L6_N0),
	.RST(SYNC_SCAN_RST1),
	.WrEn(WrEn),
	.RdEn(RdEn),
	.Address({ Address[3],
		Address[2],
		n4,
		n3 }),
	.WrData({ Wr_D[7],
		Wr_D[6],
		Wr_D[5],
		Wr_D[4],
		Wr_D[3],
		Wr_D[2],
		Wr_D[1],
		Wr_D[0] }),
	.RdData({ Rd_D[7],
		Rd_D[6],
		Rd_D[5],
		Rd_D[4],
		Rd_D[3],
		Rd_D[2],
		Rd_D[1],
		Rd_D[0] }),
	.RdData_VLD(RD_D_VLD),
	.REG0({ Op_A[7],
		Op_A[6],
		Op_A[5],
		Op_A[4],
		Op_A[3],
		Op_A[2],
		Op_A[1],
		Op_A[0] }),
	.REG1({ Op_B[7],
		Op_B[6],
		Op_B[5],
		Op_B[4],
		Op_B[3],
		Op_B[2],
		Op_B[1],
		Op_B[0] }),
	.REG2({ UART_CONFIG[7],
		UART_CONFIG[6],
		UART_CONFIG[5],
		UART_CONFIG[4],
		UART_CONFIG[3],
		UART_CONFIG[2],
		UART_CONFIG[1],
		UART_CONFIG[0] }),
	.REG3({ div_ratio[7],
		div_ratio[6],
		div_ratio[5],
		div_ratio[4],
		div_ratio[3],
		div_ratio[2],
		div_ratio[1],
		div_ratio[0] }),
	.test_si3(SI[0]),
	.test_si2(SI[1]),
	.test_si1(n15),
	.test_so2(n11),
	.test_so1(SO[1]),
	.test_se(SE),
	.FE_OFN0_SYNC_SCAN_RST1(FE_OFN0_SYNC_SCAN_RST1),
	.FE_OFN1_SYNC_SCAN_RST1(FE_OFN1_SYNC_SCAN_RST1),
	.REF_SCAN_CLK__L6_N1(REF_SCAN_CLK__L6_N1),
	.REF_SCAN_CLK__L6_N10(REF_SCAN_CLK__L6_N10),
	.REF_SCAN_CLK__L6_N11(REF_SCAN_CLK__L6_N11),
	.REF_SCAN_CLK__L6_N2(REF_SCAN_CLK__L6_N2),
	.REF_SCAN_CLK__L6_N3(REF_SCAN_CLK__L6_N3),
	.REF_SCAN_CLK__L6_N7(REF_SCAN_CLK__L6_N7),
	.REF_SCAN_CLK__L6_N8(REF_SCAN_CLK__L6_N8),
	.REF_SCAN_CLK__L6_N9(REF_SCAN_CLK__L6_N9), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_OPER_WIDTH8_test_1 ALU_INST (
	.A({ Op_A[7],
		Op_A[6],
		Op_A[5],
		Op_A[4],
		Op_A[3],
		Op_A[2],
		Op_A[1],
		Op_A[0] }),
	.B({ Op_B[7],
		Op_B[6],
		Op_B[5],
		Op_B[4],
		Op_B[3],
		Op_B[2],
		Op_B[1],
		Op_B[0] }),
	.ALU_FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }),
	.ALU_CLK(CLK_ALU__L3_N0),
	.RST(FE_OFN1_SYNC_SCAN_RST1),
	.EN(ALU_EN),
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }),
	.OUT_VALID(ALU_OUT_VLD),
	.test_si(SI[3]),
	.test_se(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   CLK_GATE CLK_GATE_INST (
	.CLK_EN(_1_net_),
	.CLK(REF_SCAN_CLK__L4_N0),
	.GATED_CLK(CLK_ALU), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M U17 (
	.Y(SO[0]),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M U18 (
	.Y(UART_TX_O),
	.A(n36), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

